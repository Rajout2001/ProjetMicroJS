-- code generated from the following source code:
--   ../vm/fail.ecl
--   ../vm/value.ecl
--   ../vm/ram.ecl
--   ../vm/frames.ecl
--   ../vm/vm.ecl
--   ../vm/main.ecl
--
-- with the following command:
--
--    ./eclat -arg=true -relax -notyB ../vm/fail.ecl ../vm/value.ecl ../vm/ram.ecl ../vm/frames.ecl ../vm/vm.ecl ../vm/main.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal run    : in std_logic;
       signal rdy    : out value(0 to 0);
       signal argument : in value(0 to 0);
       signal result : out value(0 to 0));
       
end entity;
architecture rtl of main is

  type t_state is (compute969, \$37_forever264927\, \$37_forever264928\, \$37_forever264929\, \$37_forever264930\, \$37_forever264931\, add262, copy_args_to_heap257, div259, mul260, pause_getI1000, pause_getI1008, pause_getI974, pause_getI984, pause_getI992, pause_getII1001, pause_getII1009, pause_getII975, pause_getII985, pause_getII993, pause_setI970, pause_setII971, pow258, q_wait1002, q_wait1010, q_wait972, q_wait976, q_wait986, q_wait994, sub261);
  signal \state\: t_state;
  type t_state_var1463 is (compute1281, \$105_copy_args_to_heap257\, \$106_pow258\, \$107_div259\, \$108_mul260\, \$109_sub261\, \$110_add262\, \$159_forever264955\, \$187_forever264955\, \$214_forever264955\, \$226_forever264955\, \$37_forever264955\, \$37_forever264957\, \$37_forever264958\, \$37_forever264959\, \$37_forever264960\, \$37_forever264961\, pause_getI1286, pause_getI1296, pause_getI1304, pause_getI1312, pause_getI1320, pause_getII1287, pause_getII1297, pause_getII1305, pause_getII1313, pause_getII1321, pause_setI1282, pause_setI1326, pause_setI1331, pause_setI1336, pause_setI1341, pause_setI1346, pause_setI1353, pause_setI1359, pause_setI1364, pause_setI1369, pause_setI1374, pause_setI1381, pause_setI1387, pause_setI1392, pause_setI1397, pause_setI1402, pause_setI1409, pause_setI1414, pause_setI1419, pause_setI1424, pause_setI1430, pause_setI1435, pause_setI1440, pause_setI1446, pause_setI1451, pause_setII1283, pause_setII1327, pause_setII1332, pause_setII1337, pause_setII1342, pause_setII1347, pause_setII1354, pause_setII1360, pause_setII1365, pause_setII1370, pause_setII1375, pause_setII1382, pause_setII1388, pause_setII1393, pause_setII1398, pause_setII1403, pause_setII1410, pause_setII1415, pause_setII1420, pause_setII1425, pause_setII1431, pause_setII1436, pause_setII1441, pause_setII1447, pause_setII1452, q_wait1284, q_wait1288, q_wait1298, q_wait1306, q_wait1314, q_wait1322, q_wait1328, q_wait1333, q_wait1338, q_wait1343, q_wait1348, q_wait1355, q_wait1361, q_wait1366, q_wait1371, q_wait1376, q_wait1383, q_wait1389, q_wait1394, q_wait1399, q_wait1404, q_wait1411, q_wait1416, q_wait1421, q_wait1426, q_wait1432, q_wait1437, q_wait1442, q_wait1448, q_wait1453);
  signal state_var1463: t_state_var1463;
  type t_state_var1462 is (compute1278);
  signal state_var1462: t_state_var1462;
  type t_state_var1461 is (compute1273);
  signal state_var1461: t_state_var1461;
  type t_state_var1460 is (compute1016, \$37_forever264932\, \$37_forever264934\, \$37_forever264935\, \$37_forever264936\, \$37_forever264937\, \$37_forever264938\, \$37_forever264944\, \$37_forever264945\, \$37_forever264946\, \$37_forever264947\, \$37_forever264948\, \$37_forever264949\, \$37_forever264950\, \$37_forever264951\, \$37_forever264952\, \$37_forever264953\, \$37_forever264954\, \$39_copy_args_to_heap257\, \$40_pow258\, \$41_div259\, \$42_mul260\, \$43_sub261\, \$44_add262\, \$63_forever264932\, \$76_forever264932\, \$87_forever264932\, \$95_forever264932\, forever263933, forever263939, forever263940, forever263941, forever263942, forever263943, pause_getI1021, pause_getI1031, pause_getI1039, pause_getI1047, pause_getI1055, pause_getI1093, pause_getI1097, pause_getI1110, pause_getI1117, pause_getI1129, pause_getI1136, pause_getI1148, pause_getI1165, pause_getI1178, pause_getI1185, pause_getI1192, pause_getI1200, pause_getI1213, pause_getI1217, pause_getI1225, pause_getI1236, pause_getI1249, pause_getI1257, pause_getI1263, pause_getII1022, pause_getII1032, pause_getII1040, pause_getII1048, pause_getII1056, pause_getII1094, pause_getII1098, pause_getII1111, pause_getII1118, pause_getII1130, pause_getII1137, pause_getII1149, pause_getII1166, pause_getII1179, pause_getII1186, pause_getII1193, pause_getII1201, pause_getII1214, pause_getII1218, pause_getII1226, pause_getII1237, pause_getII1250, pause_getII1258, pause_getII1264, pause_setI1017, pause_setI1063, pause_setI1067, pause_setI1072, pause_setI1077, pause_setI1103, pause_setI1122, pause_setI1141, pause_setI1153, pause_setI1158, pause_setI1170, pause_setI1196, pause_setI1205, pause_setI1209, pause_setI1221, pause_setI1241, pause_setI1245, pause_setI1253, pause_setII1018, pause_setII1064, pause_setII1068, pause_setII1073, pause_setII1078, pause_setII1104, pause_setII1123, pause_setII1142, pause_setII1154, pause_setII1159, pause_setII1171, pause_setII1197, pause_setII1206, pause_setII1210, pause_setII1222, pause_setII1242, pause_setII1246, pause_setII1254, q_wait1019, q_wait1023, q_wait1033, q_wait1041, q_wait1049, q_wait1057, q_wait1065, q_wait1069, q_wait1074, q_wait1079, q_wait1095, q_wait1099, q_wait1105, q_wait1112, q_wait1119, q_wait1124, q_wait1131, q_wait1138, q_wait1143, q_wait1150, q_wait1155, q_wait1160, q_wait1167, q_wait1172, q_wait1180, q_wait1187, q_wait1194, q_wait1198, q_wait1202, q_wait1207, q_wait1211, q_wait1215, q_wait1219, q_wait1223, q_wait1227, q_wait1238, q_wait1243, q_wait1247, q_wait1251, q_wait1255, q_wait1259, q_wait1265, vm_run_code247);
  signal state_var1460: t_state_var1460;
  type array_value_68 is array (natural range <>) of value(0 to 67);
  type array_value_72 is array (natural range <>) of value(0 to 71);
  type array_value_128 is array (natural range <>) of value(0 to 127);
  signal arr962 : array_value_68(0 to 99) := (others => (others => '0'));
  signal \$arr962_value\ : value(0 to 67);
  signal \$arr962_ptr\ : natural range 0 to 99;
  signal \$arr962_ptr_write\ : natural range 0 to 99;
  signal \$arr962_write\ : value(0 to 67);
  signal \$arr962_write_request\ : std_logic := '0';
  signal arr963 : array_value_68(0 to 99) := (others => (others => '0'));
  signal \$arr963_value\ : value(0 to 67);
  signal \$arr963_ptr\ : natural range 0 to 99;
  signal \$arr963_ptr_write\ : natural range 0 to 99;
  signal \$arr963_write\ : value(0 to 67);
  signal \$arr963_write_request\ : std_logic := '0';
  signal arr964 : array_value_68(0 to 99) := (others => (others => '0'));
  signal \$arr964_value\ : value(0 to 67);
  signal \$arr964_ptr\ : natural range 0 to 99;
  signal \$arr964_ptr_write\ : natural range 0 to 99;
  signal \$arr964_write\ : value(0 to 67);
  signal \$arr964_write_request\ : std_logic := '0';
  signal arr965 : array_value_72(0 to 99) := (others => (others => '0'));
  signal \$arr965_value\ : value(0 to 71);
  signal \$arr965_ptr\ : natural range 0 to 99;
  signal \$arr965_ptr_write\ : natural range 0 to 99;
  signal \$arr965_write\ : value(0 to 71);
  signal \$arr965_write_request\ : std_logic := '0';
  signal arr966 : array_value_128(0 to 99) := (others => (others => '0'));
  signal \$arr966_value\ : value(0 to 127);
  signal \$arr966_ptr\ : natural range 0 to 99;
  signal \$arr966_ptr_write\ : natural range 0 to 99;
  signal \$arr966_write\ : value(0 to 127);
  signal \$arr966_write_request\ : std_logic := '0';
  
  begin
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr962_write_request\ = '1' then
                    arr962(\$arr962_ptr_write\) <= \$arr962_write\;
                  else
                   \$arr962_value\ <= arr962(\$arr962_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr963_write_request\ = '1' then
                    arr963(\$arr963_ptr_write\) <= \$arr963_write\;
                  else
                   \$arr963_value\ <= arr963(\$arr963_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr964_write_request\ = '1' then
                    arr964(\$arr964_ptr_write\) <= \$arr964_write\;
                  else
                   \$arr964_value\ <= arr964(\$arr964_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr965_write_request\ = '1' then
                    arr965(\$arr965_ptr_write\) <= \$arr965_write\;
                  else
                   \$arr965_value\ <= arr965(\$arr965_ptr\);
                  end if;
            end if;
        end process;
    
    process (clk)
            begin
            if (rising_edge(clk)) then
                  if \$arr966_write_request\ = '1' then
                    arr966(\$arr966_ptr_write\) <= \$arr966_write\;
                  else
                   \$arr966_value\ <= arr966(\$arr966_ptr\);
                  end if;
            end if;
        end process;
    
    process(clk)
      variable \$v723\, \$v711\ : value(0 to 1) := (others => '0');
      variable mul260_arg, pow258_arg, \$44_add262_arg\, \$110_add262_arg\, 
               \$107_div259_arg\, \$109_sub261_arg\, sub261_arg, add262_arg, 
               div259_arg, \$43_sub261_arg\, \$41_div259_arg\, 
               \$106_pow258_arg\, \$108_mul260_arg\, \$42_mul260_arg\, 
               \$40_pow258_arg\ : value(0 to 95) := (others => '0');
      variable \$v1317\, \$v1189\, \$v989\, \$v1052\, \$v1036\, \$v1309\, 
               \$v1082\, \$v1088\, \$v1133\, \$v1062\, \$v1114\, \$v1145\, 
               \$v1204\, \$v1044\, \$v1162\, \$v1028\, \$v1229\, \$v1107\, 
               \$v997\, \$v1085\, \$v760\, \$v1293\, \$v1081\, \$v1005\, 
               \$v1301\, \$v1126\, \$v1182\, \$v981\ : value(0 to 63) := (others => '0');
      variable \$v1261\, instr : value(0 to 71) := (others => '0');
      variable \$39_copy_args_to_heap257_arg\, copy_args_to_heap257_arg, 
               \$105_copy_args_to_heap257_arg\ : value(0 to 159) := (others => '0');
      variable \$v1407\, \$v1231\, \$v1174\, \$v1379\, p, \$v1351\ : value(0 to 4) := (others => '0');
      variable \$v1319\, \$v1090\, \$v1128\, \$v1092\, \$v1232\, \$v1311\, 
               \$v1191\, \$v1109\, \$v991\, \$v1046\, \$v1038\, \$v1084\, 
               \$v1175\, \$v1030\, \$v1184\, \$v1007\, \$v1054\, \$v1164\, 
               \$v1295\, \$v1147\, \$v1135\, \$v1177\, \$v1303\, \$v1087\, 
               \$v1235\, \$v983\, \$v1262\, \$v999\, \$v1116\ : value(0 to 3) := (others => '0');
      variable vm_run_code247_arg : value(0 to 294) := (others => '0');
      variable \$v843\ : value(0 to 127) := (others => '0');
      variable \$v1020\, \$v1139\, \$v1454\, \$v1173\, \$v1433\, \$v1239\, 
               \$v1012\, \$v1334\, \$v1434\, \$v1216\, \$v1080\, \$v1325\, 
               \$v1324\, \$v1438\, \$v1299\, rdy1015, \$v1329\, \$v1267\, 
               \$v1362\, \$v1356\, \$v1025\, \$v1058\, result967, \$v1270\, 
               \$v1208\, \$v1443\, \$v1307\, \$v1248\, \$v1349\, \$v722\, 
               \$v1199\, \$v1027\, x, \$v1113\, \$v980\, \$34_b\, \$v1323\, 
               \$v1350\, \$v1106\, \$v1195\, \$v1125\, \$v1042\, rdy1272, 
               \$v1427\, \$v988\, \$v1100\, \$v1367\, \$v1339\, \$v1316\, 
               \$v1244\, jfalse, result1279, \$v1096\, \$v1102\, \$v1224\, 
               \$v1059\, \$v978\, \$v1075\, a1, \$v1024\, \$v1003\, \$v1291\, 
               \$v1459\, \$v1260\, \$v1315\, \$v1372\, \$v1140\, \$v1076\, 
               is_loaded, \$v1300\, \$v1308\, \$v977\, vm_run_code247_result, 
               \$v987\, \$v1051\, \$v1240\, \$v1417\, \$v1169\, \$v1252\, 
               \$v1203\, \$v1289\, b2, \$v1035\, \$v996\, \$v1457\, \$v995\, 
               \$v1228\, \$v1422\, \$v1395\, \$v1132\, result1014, \$v1026\, 
               \$v1004\, \$v1011\, \$v1292\, \$v1400\, \$v1066\, \$v1101\, 
               \$v1120\, \$v1456\, \$v1212\, \$v1290\, \$v1266\, \$v1152\, 
               \$v1390\, \$v1188\, \$v979\, \$v1050\, rdy1277, \$v1230\, 
               \$v1256\, \$v1121\, rdy968, \$v1233\, \$v1377\, \$v1378\, 
               \$v1156\, \$v1070\, \$v1144\, \$v1268\, \$v1161\, \$v1405\, 
               \$v1406\, \$v1181\, \$v1344\, \$v1013\, \$v973\, rdy1280, 
               \$v1151\, \$v1060\, \$v1043\, verif, \$v1220\, \$v1384\, 
               \$v1450\, \$v1412\, \$v1275\, result1276, \$v1285\, \$v1449\, 
               jtrue, \$v1034\, \$v1168\ : value(0 to 0) := (others => '0');
      variable \$325_a\, \$v1357\, \$40_pow258_result\, \$v1373\, i, 
               \$41_div259_result\, \$v1439\, \$59_a\, \$v1444\, \$20_l\, 
               \$v1363\, \$356_a\, cy, puissance, addition, mult, 
               \$296_sous\, \$v1368\, divisor, l, 
               \$39_copy_args_to_heap257_result\, \$v1401\, \$91_a\, sous, 
               \$21_i\, \$v721\, \$17_l\, n, \$44_add262_result\, res, 
               \$v1385\, \$v1428\, \$v1345\, \$v1335\, \$v1391\, 
               \$343_divisor\, \$19_i\, \$33_n\, \$202_divisor\, \$v1340\, 
               \$72_a\, \$147_sous\, \$180_a\, valeur_depart, \$175_mult\, 
               \$320_mult\, \$v1157\, \$125_a\, \$120_addition\, \$18_l\, 
               \$22_i\, \$v1396\, \$v1330\, resultat, \$v1423\, \$v1071\, 
               result1271, \$301_a\, \$v1418\, \$277_a\, b, \$152_a\, 
               \$43_sub261_result\, \$219_a\, \$272_addition\, 
               \$42_mul260_result\, \$v1413\, a : value(0 to 31) := (others => '0');
      variable \$v752\ : value(0 to 293) := (others => '0');
      variable \$v1045\, \$v1352\, \$271_var\, \$259\, \$71_var\, \$v1115\, 
               \$v111\, \$v990\, \$v1445\, \$v1061\, \$v1108\, \$319_var\, 
               temp, \$v982\, \$v52\, \$v1294\, \$v1310\, \$v1183\, \$v165\, 
               \$295_var\, \$v13\, \$v1127\, \$58_var\, e1, \$v170\, 
               \$v1146\, \$v1006\, \$v1234\, \$v1386\, \$v43\, var, \$v1037\, 
               \$v1134\, \$v1083\, \$218\, e2, \$v1190\, \$v1358\, \$v1029\, 
               \$392\, \$v41\, \$v151\, \$v998\, \$146_var\, \$v1086\, 
               \value\, \$v174\, \$v70\, \$v1429\, \$v1176\, \$v78\, 
               \$v1318\, \$355\, \$119_var\, \$v54\, \$v1302\, \$v1408\, 
               \$v1053\, \$v1089\, \$v1091\, \$174_var\, v, \$v1163\, 
               \$v1380\ : value(0 to 67) := (others => '0');
      variable \$arr962_ptr_take\ : value(0 to 0) := "0";
      variable \$arr963_ptr_take\ : value(0 to 0) := "0";
      variable \$arr964_ptr_take\ : value(0 to 0) := "0";
      variable \$arr965_ptr_take\ : value(0 to 0) := "0";
      variable \$arr966_ptr_take\ : value(0 to 0) := "0";
      
    begin
      
      if rising_edge(clk) then
        if (reset = '1') then
          default_zero(a); default_zero(\$v1380\); default_zero(\$v1116\); 
          default_zero(\$v981\); default_zero(\$v1168\); 
          default_zero(\$v1351\); default_zero(\$v1034\); 
          default_zero(\$v1163\); default_zero(\$v1182\); 
          default_zero(\$v1413\); default_zero(jtrue); 
          default_zero(\$42_mul260_result\); default_zero(\$40_pow258_arg\); 
          default_zero(\$v1449\); default_zero(\$v1285\); 
          default_zero(\$v999\); default_zero(v); default_zero(\$v711\); 
          default_zero(result1276); default_zero(\$272_addition\); 
          default_zero(\$219_a\); default_zero(\$v1275\); 
          default_zero(\$v1412\); default_zero(\$42_mul260_arg\); 
          default_zero(\$v1262\); default_zero(\$174_var\); 
          default_zero(\$v1450\); default_zero(\$43_sub261_result\); 
          default_zero(\$152_a\); default_zero(\$v1091\); 
          default_zero(\$v1089\); default_zero(b); default_zero(\$v1384\); 
          default_zero(\$v1220\); default_zero(verif); 
          default_zero(\$v1043\); default_zero(\$277_a\); 
          default_zero(\$v1053\); default_zero(vm_run_code247_arg); 
          default_zero(\$v1418\); default_zero(\$301_a\); 
          default_zero(\$v1060\); default_zero(\$v1126\); 
          default_zero(\$v983\); default_zero(\$v1151\); 
          default_zero(\$v1301\); default_zero(rdy1280); 
          default_zero(\$v973\); default_zero(\$108_mul260_arg\); 
          default_zero(\$v1013\); default_zero(\$v1408\); 
          default_zero(\$v1344\); default_zero(\$v1005\); 
          default_zero(\$v1181\); default_zero(\$v1406\); 
          default_zero(\$v1405\); default_zero(\$v1302\); 
          default_zero(\$v1081\); default_zero(\$v1161\); 
          default_zero(result1271); default_zero(\$106_pow258_arg\); 
          default_zero(\$v1268\); default_zero(\$v1235\); 
          default_zero(\$v1144\); default_zero(\$v1087\); 
          default_zero(\$v1070\); default_zero(\$v1303\); 
          default_zero(\$v1071\); default_zero(\$v1156\); 
          default_zero(\$v1378\); default_zero(\$v1423\); 
          default_zero(\$v1377\); default_zero(\$v54\); 
          default_zero(\$v1233\); default_zero(\$v1177\); 
          default_zero(resultat); default_zero(rdy968); 
          default_zero(\$v1121\); default_zero(\$41_div259_arg\); 
          default_zero(\$119_var\); default_zero(\$v1256\); 
          default_zero(\$355\); default_zero(\$v1318\); 
          default_zero(\$v1230\); default_zero(\$v1330\); 
          default_zero(rdy1277); default_zero(\$v1135\); 
          default_zero(\$43_sub261_arg\); default_zero(\$v78\); 
          default_zero(\$v1050\); default_zero(\$v843\); 
          default_zero(\$v1147\); default_zero(\$v979\); 
          default_zero(\$v1188\); default_zero(\$v1176\); 
          default_zero(\$v1295\); default_zero(\$v1396\); 
          default_zero(\$v1429\); default_zero(\$v1390\); 
          default_zero(\$v1152\); default_zero(\$v70\); 
          default_zero(\$v1266\); default_zero(\$v1293\); 
          default_zero(\$v1290\); default_zero(\$v174\); 
          default_zero(\$v1212\); default_zero(div259_arg); 
          default_zero(\$v1456\); default_zero(add262_arg); default_zero(p); 
          default_zero(\value\); default_zero(\$v1120\); 
          default_zero(\$v1086\); default_zero(\$v1101\); 
          default_zero(\$v1066\); default_zero(\$22_i\); 
          default_zero(\$v1164\); default_zero(\$v760\); 
          default_zero(\$v1400\); default_zero(\$146_var\); 
          default_zero(\$v1292\); default_zero(\$v1011\); 
          default_zero(\$v1004\); default_zero(sub261_arg); 
          default_zero(\$v1026\); default_zero(result1014); 
          default_zero(\$18_l\); default_zero(\$v1132\); 
          default_zero(\$120_addition\); default_zero(\$v1395\); 
          default_zero(\$v1422\); default_zero(\$v998\); 
          default_zero(\$v1228\); default_zero(\$v1085\); 
          default_zero(\$125_a\); default_zero(\$v995\); 
          default_zero(\$v1157\); default_zero(\$v1457\); 
          default_zero(\$v1054\); default_zero(\$v1379\); 
          default_zero(\$v996\); default_zero(\$v1035\); 
          default_zero(\$109_sub261_arg\); default_zero(\$v151\); 
          default_zero(b2); default_zero(\$v41\); default_zero(\$320_mult\); 
          default_zero(\$v723\); default_zero(\$392\); 
          default_zero(\$v1289\); default_zero(\$v1029\); 
          default_zero(\$v1358\); default_zero(\$v1007\); 
          default_zero(\$v1190\); default_zero(\$175_mult\); 
          default_zero(valeur_depart); default_zero(\$v1203\); 
          default_zero(e2); default_zero(\$218\); default_zero(\$v997\); 
          default_zero(\$v1252\); default_zero(\$v1083\); 
          default_zero(\$v1169\); default_zero(\$v1417\); 
          default_zero(\$v1240\); default_zero(\$180_a\); 
          default_zero(\$v1174\); default_zero(\$v1107\); 
          default_zero(\$147_sous\); default_zero(\$v1229\); 
          default_zero(\$v1051\); default_zero(\$72_a\); 
          default_zero(\$v1184\); default_zero(\$v987\); 
          default_zero(\$v1028\); default_zero(\$v1340\); 
          default_zero(\$202_divisor\); default_zero(vm_run_code247_result); 
          default_zero(\$v1134\); default_zero(\$v1037\); 
          default_zero(\$v977\); 
          default_zero(\$105_copy_args_to_heap257_arg\); 
          default_zero(\$33_n\); default_zero(var); default_zero(\$v1308\); 
          default_zero(\$v1300\); default_zero(is_loaded); 
          default_zero(\$v1076\); default_zero(\$19_i\); 
          default_zero(\$v1140\); default_zero(copy_args_to_heap257_arg); 
          default_zero(\$343_divisor\); default_zero(\$v1030\); 
          default_zero(\$v752\); default_zero(\$v1162\); 
          default_zero(\$v1391\); default_zero(\$v1372\); 
          default_zero(\$v1335\); default_zero(\$v1315\); 
          default_zero(\$v1260\); default_zero(\$v1345\); 
          default_zero(\$v1459\); default_zero(\$v1291\); 
          default_zero(\$v1428\); default_zero(\$107_div259_arg\); 
          default_zero(\$v43\); default_zero(\$v1044\); 
          default_zero(\$v1003\); default_zero(\$v1024\); 
          default_zero(\$v1175\); default_zero(a1); default_zero(\$v1385\); 
          default_zero(res); default_zero(\$v1075\); default_zero(\$v1084\); 
          default_zero(\$v1204\); default_zero(\$44_add262_result\); 
          default_zero(\$v1386\); default_zero(\$v978\); 
          default_zero(\$v1059\); default_zero(\$v1224\); 
          default_zero(\$v1102\); default_zero(n); default_zero(\$v1231\); 
          default_zero(\$17_l\); default_zero(\$v1096\); 
          default_zero(result1279); default_zero(jfalse); 
          default_zero(\$v1244\); default_zero(\$v721\); 
          default_zero(\$v1316\); default_zero(\$v1339\); 
          default_zero(\$v1145\); default_zero(\$v1367\); 
          default_zero(\$v1100\); default_zero(\$v1114\); 
          default_zero(\$v1062\); default_zero(\$21_i\); 
          default_zero(\$v988\); default_zero(\$v1234\); 
          default_zero(\$v1427\); default_zero(sous); default_zero(rdy1272); 
          default_zero(\$v1006\); default_zero(\$91_a\); 
          default_zero(\$v1133\); default_zero(\$v1401\); 
          default_zero(\$v1042\); default_zero(\$v1146\); 
          default_zero(\$v1125\); 
          default_zero(\$39_copy_args_to_heap257_result\); 
          default_zero(\$v1195\); default_zero(\$v170\); 
          default_zero(\$v1038\); default_zero(e1); default_zero(l); 
          default_zero(\$v1106\); default_zero(\$58_var\); 
          default_zero(\$v1046\); default_zero(\$v1350\); 
          default_zero(instr); default_zero(\$v1088\); default_zero(divisor); 
          default_zero(\$v1127\); default_zero(\$v13\); 
          default_zero(\$v1323\); default_zero(\$34_b\); 
          default_zero(\$v1368\); default_zero(\$295_var\); 
          default_zero(\$296_sous\); default_zero(\$v165\); 
          default_zero(\$v980\); default_zero(\$v1183\); 
          default_zero(\$v1082\); default_zero(\$v1309\); 
          default_zero(\$v1310\); default_zero(\$v991\); 
          default_zero(\$v1113\); default_zero(x); default_zero(\$v1294\); 
          default_zero(mult); default_zero(\$v1036\); default_zero(\$v1027\); 
          default_zero(addition); default_zero(\$v1199\); 
          default_zero(puissance); default_zero(\$110_add262_arg\); 
          default_zero(\$v52\); default_zero(\$v722\); default_zero(cy); 
          default_zero(\$v1349\); default_zero(\$v982\); 
          default_zero(\$v1248\); default_zero(\$v1109\); 
          default_zero(\$v1307\); default_zero(\$356_a\); 
          default_zero(\$v1443\); default_zero(\$v1363\); 
          default_zero(\$v1208\); default_zero(temp); default_zero(\$v1270\); 
          default_zero(\$v1407\); default_zero(result967); 
          default_zero(\$20_l\); default_zero(\$v1444\); 
          default_zero(\$v1058\); default_zero(\$v1025\); 
          default_zero(\$319_var\); default_zero(\$59_a\); 
          default_zero(\$v1356\); default_zero(\$v1362\); 
          default_zero(\$v1439\); default_zero(\$v1108\); 
          default_zero(\$v1267\); default_zero(\$v1329\); 
          default_zero(rdy1015); default_zero(\$44_add262_arg\); 
          default_zero(\$v1299\); default_zero(\$v1052\); 
          default_zero(\$41_div259_result\); default_zero(\$v1261\); 
          default_zero(i); default_zero(\$v1438\); default_zero(\$v1061\); 
          default_zero(\$39_copy_args_to_heap257_arg\); 
          default_zero(\$v1445\); default_zero(\$v1324\); 
          default_zero(\$v1373\); default_zero(\$v990\); 
          default_zero(\$v1191\); default_zero(\$40_pow258_result\); 
          default_zero(\$v1325\); default_zero(\$v1357\); 
          default_zero(\$v989\); default_zero(\$v1080\); 
          default_zero(\$325_a\); default_zero(\$v111\); 
          default_zero(\$v1216\); default_zero(\$v1434\); 
          default_zero(\$v1115\); default_zero(\$v1334\); 
          default_zero(\$v1012\); default_zero(\$v1311\); 
          default_zero(\$71_var\); default_zero(\$v1239\); 
          default_zero(\$v1232\); default_zero(\$v1189\); 
          default_zero(\$259\); default_zero(\$v1433\); 
          default_zero(\$v1092\); default_zero(\$v1173\); 
          default_zero(\$271_var\); default_zero(\$v1454\); 
          default_zero(\$v1139\); default_zero(pow258_arg); 
          default_zero(\$v1317\); default_zero(mul260_arg); 
          default_zero(\$v1352\); default_zero(\$v1128\); 
          default_zero(\$v1090\); default_zero(\$v1319\); 
          default_zero(\$v1045\); default_zero(\$v1020\); 
          rdy <= "1";
          rdy968 := "0";
          \state\ <= compute969;
          state_var1463 <= compute1281;
          state_var1462 <= compute1278;
          state_var1461 <= compute1273;
          state_var1460 <= compute1016;
          
        else if run = '1' then
          case \state\ is
          when \$37_forever264927\ =>
            \state\ <= \$37_forever264927\;
          when \$37_forever264928\ =>
            \state\ <= \$37_forever264928\;
          when \$37_forever264929\ =>
            \state\ <= \$37_forever264929\;
          when \$37_forever264930\ =>
            \state\ <= \$37_forever264930\;
          when \$37_forever264931\ =>
            \state\ <= \$37_forever264931\;
          when add262 =>
            \$v1012\ := eclat_eq(add262_arg(0 to 31) & "00000000000000000000000000000000");
            if \$v1012\(0) = '1' then
              \state\ <= add262;
            else
              \$v1011\ := \$arr963_ptr_take\;
              if \$v1011\(0) = '1' then
                \state\ <= q_wait1010;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(add262_arg(64 to 95) & "00000000000000000000000000000001") & add262_arg(0 to 31))));
                \state\ <= pause_getI1008;
              end if;
            end if;
          when copy_args_to_heap257 =>
            \$v978\ := eclat_eq(copy_args_to_heap257_arg(0 to 31) & "00000000000000000000000000000000");
            if \$v978\(0) = '1' then
              \state\ <= copy_args_to_heap257;
            else
              \$v977\ := \$arr963_ptr_take\;
              if \$v977\(0) = '1' then
                \state\ <= q_wait976;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(copy_args_to_heap257_arg(96 to 127) & copy_args_to_heap257_arg(0 to 31)) & "00000000000000000000000000000001")));
                \state\ <= pause_getI974;
              end if;
            end if;
          when div259 =>
            \$v988\ := eclat_eq(div259_arg(0 to 31) & "00000000000000000000000000000000");
            if \$v988\(0) = '1' then
              \state\ <= div259;
            else
              \$v987\ := \$arr963_ptr_take\;
              if \$v987\(0) = '1' then
                \state\ <= q_wait986;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(div259_arg(64 to 95) & "00000000000000000000000000000001") & div259_arg(0 to 31))));
                \state\ <= pause_getI984;
              end if;
            end if;
          when mul260 =>
            \$v996\ := eclat_eq(mul260_arg(0 to 31) & "00000000000000000000000000000000");
            if \$v996\(0) = '1' then
              \state\ <= mul260;
            else
              \$v995\ := \$arr963_ptr_take\;
              if \$v995\(0) = '1' then
                \state\ <= q_wait994;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(mul260_arg(64 to 95) & "00000000000000000000000000000001") & mul260_arg(0 to 31))));
                \state\ <= pause_getI992;
              end if;
            end if;
          when pause_getI1000 =>
            \state\ <= pause_getII1001;
          when pause_getI1008 =>
            \state\ <= pause_getII1009;
          when pause_getI974 =>
            \state\ <= pause_getII975;
          when pause_getI984 =>
            \state\ <= pause_getII985;
          when pause_getI992 =>
            \state\ <= pause_getII993;
          when pause_getII1001 =>
            \$arr963_ptr_take\(0) := '0';
            \$295_var\ := \$arr963_value\;
            \$v998\ := \$295_var\;
            \$v999\ := \$v998\(0 to 3);
            \$v997\ := \$v998\(4 to 67);
            case \$v999\ is
            when "0001" =>
              \$301_a\ := \$v997\(0 to 31);
              \$296_sous\ := \$301_a\;
              sub261_arg := eclat_sub(sub261_arg(0 to 31) & "00000000000000000000000000000001") & eclat_sub(sub261_arg(32 to 63) & \$296_sous\) & sub261_arg(64 to 95);
              \state\ <= sub261;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("NON INT"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$37_forever264930\;
            end case;
          when pause_getII1009 =>
            \$arr963_ptr_take\(0) := '0';
            \$271_var\ := \$arr963_value\;
            \$v1006\ := \$271_var\;
            \$v1007\ := \$v1006\(0 to 3);
            \$v1005\ := \$v1006\(4 to 67);
            case \$v1007\ is
            when "0001" =>
              \$277_a\ := \$v1005\(0 to 31);
              \$272_addition\ := \$277_a\;
              add262_arg := eclat_sub(add262_arg(0 to 31) & "00000000000000000000000000000001") & eclat_add(add262_arg(32 to 63) & \$272_addition\) & add262_arg(64 to 95);
              \state\ <= add262;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("NON INT "));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$37_forever264931\;
            end case;
          when pause_getII975 =>
            \$arr963_ptr_take\(0) := '0';
            \$392\ := \$arr963_value\;
            \$v973\ := \$arr962_ptr_take\;
            if \$v973\(0) = '1' then
              \state\ <= q_wait972;
            else
              \$arr962_ptr_take\(0) := '1';
              \$arr962_ptr_write\ <= to_integer(unsigned(copy_args_to_heap257_arg(128 to 159)));
              \$arr962_write_request\ <= '1';
              \$arr962_write\ <= \$392\;
              \state\ <= pause_setI970;
            end if;
          when pause_getII985 =>
            \$arr963_ptr_take\(0) := '0';
            \$355\ := \$arr963_value\;
            \$v982\ := \$355\;
            \$v983\ := \$v982\(0 to 3);
            \$v981\ := \$v982\(4 to 67);
            case \$v983\ is
            when "0001" =>
              \$356_a\ := \$v981\(0 to 31);
              \$343_divisor\ := \$356_a\;
              \$v980\ := eclat_eq(\$343_divisor\ & "00000000000000000000000000000000");
              if \$v980\(0) = '1' then
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("Div par zero impossible"));
                
                eclat_print_newline(eclat_unit);
                
                \state\ <= \$37_forever264927\;
              else
                div259_arg := eclat_sub(div259_arg(0 to 31) & "00000000000000000000000000000001") & eclat_div(div259_arg(32 to 63) & \$343_divisor\) & div259_arg(64 to 95);
                \state\ <= div259;
              end if;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("NON INT"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$37_forever264928\;
            end case;
          when pause_getII993 =>
            \$arr963_ptr_take\(0) := '0';
            \$319_var\ := \$arr963_value\;
            \$v990\ := \$319_var\;
            \$v991\ := \$v990\(0 to 3);
            \$v989\ := \$v990\(4 to 67);
            case \$v991\ is
            when "0001" =>
              \$325_a\ := \$v989\(0 to 31);
              \$320_mult\ := \$325_a\;
              mul260_arg := eclat_sub(mul260_arg(0 to 31) & "00000000000000000000000000000001") & eclat_mult(mul260_arg(32 to 63) & \$320_mult\) & mul260_arg(64 to 95);
              \state\ <= mul260;
            when others =>
              eclat_print_string(of_string("fatal error: "));
              
              eclat_print_string(of_string("NON INT"));
              
              eclat_print_newline(eclat_unit);
              
              \state\ <= \$37_forever264929\;
            end case;
          when pause_setI970 =>
            \$arr962_write_request\ <= '0';
            \state\ <= pause_setII971;
          when pause_setII971 =>
            \$arr962_ptr_take\(0) := '0';
            copy_args_to_heap257_arg := eclat_sub(copy_args_to_heap257_arg(0 to 31) & "00000000000000000000000000000001") & copy_args_to_heap257_arg(32 to 63) & eclat_add(copy_args_to_heap257_arg(64 to 95) & "00000000000000000000000000000001") & copy_args_to_heap257_arg(96 to 127) & copy_args_to_heap257_arg(128 to 159);
            \state\ <= copy_args_to_heap257;
          when pow258 =>
            \$v979\ := eclat_eq(pow258_arg(32 to 63) & "00000000000000000000000000000000");
            if \$v979\(0) = '1' then
              \state\ <= pow258;
            else
              pow258_arg := pow258_arg(0 to 31) & eclat_sub(pow258_arg(32 to 63) & "00000000000000000000000000000001") & eclat_mult(pow258_arg(64 to 95) & pow258_arg(0 to 31));
              \state\ <= pow258;
            end if;
          when q_wait1002 =>
            \$v1003\ := \$arr963_ptr_take\;
            if \$v1003\(0) = '1' then
              \state\ <= q_wait1002;
            else
              \$arr963_ptr_take\(0) := '1';
              \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(sub261_arg(64 to 95) & "00000000000000000000000000000001") & sub261_arg(0 to 31))));
              \state\ <= pause_getI1000;
            end if;
          when q_wait1010 =>
            \$v1011\ := \$arr963_ptr_take\;
            if \$v1011\(0) = '1' then
              \state\ <= q_wait1010;
            else
              \$arr963_ptr_take\(0) := '1';
              \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(add262_arg(64 to 95) & "00000000000000000000000000000001") & add262_arg(0 to 31))));
              \state\ <= pause_getI1008;
            end if;
          when q_wait972 =>
            \$v973\ := \$arr962_ptr_take\;
            if \$v973\(0) = '1' then
              \state\ <= q_wait972;
            else
              \$arr962_ptr_take\(0) := '1';
              \$arr962_ptr_write\ <= to_integer(unsigned(copy_args_to_heap257_arg(128 to 159)));
              \$arr962_write_request\ <= '1';
              \$arr962_write\ <= \$392\;
              \state\ <= pause_setI970;
            end if;
          when q_wait976 =>
            \$v977\ := \$arr963_ptr_take\;
            if \$v977\(0) = '1' then
              \state\ <= q_wait976;
            else
              \$arr963_ptr_take\(0) := '1';
              \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(copy_args_to_heap257_arg(96 to 127) & copy_args_to_heap257_arg(0 to 31)) & "00000000000000000000000000000001")));
              \state\ <= pause_getI974;
            end if;
          when q_wait986 =>
            \$v987\ := \$arr963_ptr_take\;
            if \$v987\(0) = '1' then
              \state\ <= q_wait986;
            else
              \$arr963_ptr_take\(0) := '1';
              \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(div259_arg(64 to 95) & "00000000000000000000000000000001") & div259_arg(0 to 31))));
              \state\ <= pause_getI984;
            end if;
          when q_wait994 =>
            \$v995\ := \$arr963_ptr_take\;
            if \$v995\(0) = '1' then
              \state\ <= q_wait994;
            else
              \$arr963_ptr_take\(0) := '1';
              \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(mul260_arg(64 to 95) & "00000000000000000000000000000001") & mul260_arg(0 to 31))));
              \state\ <= pause_getI992;
            end if;
          when sub261 =>
            \$v1004\ := eclat_eq(sub261_arg(0 to 31) & "00000000000000000000000000000000");
            if \$v1004\(0) = '1' then
              \state\ <= sub261;
            else
              \$v1003\ := \$arr963_ptr_take\;
              if \$v1003\(0) = '1' then
                \state\ <= q_wait1002;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(sub261_arg(64 to 95) & "00000000000000000000000000000001") & sub261_arg(0 to 31))));
                \state\ <= pause_getI1000;
              end if;
            end if;
          when compute969 =>
            rdy968 := eclat_false;
            case state_var1462 is
            when compute1278 =>
              rdy1277 := eclat_false;
              \$v1457\ := \$v722\;
              if \$v1457\(0) = '1' then
                result1276 := eclat_true;
                rdy1277 := eclat_true;
                state_var1462 <= compute1278;
              else
                case state_var1463 is
                when \$105_copy_args_to_heap257\ =>
                  \$v1290\ := eclat_eq(\$105_copy_args_to_heap257_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v1290\(0) = '1' then
                    state_var1463 <= \$105_copy_args_to_heap257\;
                  else
                    \$v1289\ := \$arr963_ptr_take\;
                    if \$v1289\(0) = '1' then
                      state_var1463 <= q_wait1288;
                    else
                      \$arr963_ptr_take\(0) := '1';
                      \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$105_copy_args_to_heap257_arg\(96 to 127) & \$105_copy_args_to_heap257_arg\(0 to 31)) & "00000000000000000000000000000001")));
                      state_var1463 <= pause_getI1286;
                    end if;
                  end if;
                when \$106_pow258\ =>
                  \$v1291\ := eclat_eq(\$106_pow258_arg\(32 to 63) & "00000000000000000000000000000000");
                  if \$v1291\(0) = '1' then
                    state_var1463 <= \$106_pow258\;
                  else
                    \$106_pow258_arg\ := \$106_pow258_arg\(0 to 31) & eclat_sub(\$106_pow258_arg\(32 to 63) & "00000000000000000000000000000001") & eclat_mult(\$106_pow258_arg\(64 to 95) & \$106_pow258_arg\(0 to 31));
                    state_var1463 <= \$106_pow258\;
                  end if;
                when \$107_div259\ =>
                  \$v1300\ := eclat_eq(\$107_div259_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v1300\(0) = '1' then
                    state_var1463 <= \$107_div259\;
                  else
                    \$v1299\ := \$arr963_ptr_take\;
                    if \$v1299\(0) = '1' then
                      state_var1463 <= q_wait1298;
                    else
                      \$arr963_ptr_take\(0) := '1';
                      \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$107_div259_arg\(64 to 95) & "00000000000000000000000000000001") & \$107_div259_arg\(0 to 31))));
                      state_var1463 <= pause_getI1296;
                    end if;
                  end if;
                when \$108_mul260\ =>
                  \$v1308\ := eclat_eq(\$108_mul260_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v1308\(0) = '1' then
                    state_var1463 <= \$108_mul260\;
                  else
                    \$v1307\ := \$arr963_ptr_take\;
                    if \$v1307\(0) = '1' then
                      state_var1463 <= q_wait1306;
                    else
                      \$arr963_ptr_take\(0) := '1';
                      \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$108_mul260_arg\(64 to 95) & "00000000000000000000000000000001") & \$108_mul260_arg\(0 to 31))));
                      state_var1463 <= pause_getI1304;
                    end if;
                  end if;
                when \$109_sub261\ =>
                  \$v1316\ := eclat_eq(\$109_sub261_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v1316\(0) = '1' then
                    state_var1463 <= \$109_sub261\;
                  else
                    \$v1315\ := \$arr963_ptr_take\;
                    if \$v1315\(0) = '1' then
                      state_var1463 <= q_wait1314;
                    else
                      \$arr963_ptr_take\(0) := '1';
                      \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$109_sub261_arg\(64 to 95) & "00000000000000000000000000000001") & \$109_sub261_arg\(0 to 31))));
                      state_var1463 <= pause_getI1312;
                    end if;
                  end if;
                when \$110_add262\ =>
                  \$v1324\ := eclat_eq(\$110_add262_arg\(0 to 31) & "00000000000000000000000000000000");
                  if \$v1324\(0) = '1' then
                    state_var1463 <= \$110_add262\;
                  else
                    \$v1323\ := \$arr963_ptr_take\;
                    if \$v1323\(0) = '1' then
                      state_var1463 <= q_wait1322;
                    else
                      \$arr963_ptr_take\(0) := '1';
                      \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$110_add262_arg\(64 to 95) & "00000000000000000000000000000001") & \$110_add262_arg\(0 to 31))));
                      state_var1463 <= pause_getI1320;
                    end if;
                  end if;
                when \$159_forever264955\ =>
                  state_var1463 <= \$159_forever264955\;
                when \$187_forever264955\ =>
                  state_var1463 <= \$187_forever264955\;
                when \$214_forever264955\ =>
                  state_var1463 <= \$214_forever264955\;
                when \$226_forever264955\ =>
                  state_var1463 <= \$226_forever264955\;
                when \$37_forever264955\ =>
                  state_var1463 <= \$37_forever264955\;
                when \$37_forever264957\ =>
                  state_var1463 <= \$214_forever264955\;
                when \$37_forever264958\ =>
                  state_var1463 <= \$226_forever264955\;
                when \$37_forever264959\ =>
                  state_var1463 <= \$187_forever264955\;
                when \$37_forever264960\ =>
                  state_var1463 <= \$159_forever264955\;
                when \$37_forever264961\ =>
                  state_var1463 <= \$37_forever264955\;
                when pause_getI1286 =>
                  state_var1463 <= pause_getII1287;
                when pause_getI1296 =>
                  state_var1463 <= pause_getII1297;
                when pause_getI1304 =>
                  state_var1463 <= pause_getII1305;
                when pause_getI1312 =>
                  state_var1463 <= pause_getII1313;
                when pause_getI1320 =>
                  state_var1463 <= pause_getII1321;
                when pause_getII1287 =>
                  \$arr963_ptr_take\(0) := '0';
                  \$259\ := \$arr963_value\;
                  \$v1285\ := \$arr962_ptr_take\;
                  if \$v1285\(0) = '1' then
                    state_var1463 <= q_wait1284;
                  else
                    \$arr962_ptr_take\(0) := '1';
                    \$arr962_ptr_write\ <= to_integer(unsigned(\$105_copy_args_to_heap257_arg\(128 to 159)));
                    \$arr962_write_request\ <= '1';
                    \$arr962_write\ <= \$259\;
                    state_var1463 <= pause_setI1282;
                  end if;
                when pause_getII1297 =>
                  \$arr963_ptr_take\(0) := '0';
                  \$218\ := \$arr963_value\;
                  \$v1294\ := \$218\;
                  \$v1295\ := \$v1294\(0 to 3);
                  \$v1293\ := \$v1294\(4 to 67);
                  case \$v1295\ is
                  when "0001" =>
                    \$219_a\ := \$v1293\(0 to 31);
                    \$202_divisor\ := \$219_a\;
                    \$v1292\ := eclat_eq(\$202_divisor\ & "00000000000000000000000000000000");
                    if \$v1292\(0) = '1' then
                      eclat_print_string(of_string("fatal error: "));
                      
                      eclat_print_string(of_string("Div par zero impossible"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      state_var1463 <= \$37_forever264957\;
                    else
                      \$107_div259_arg\ := eclat_sub(\$107_div259_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_div(\$107_div259_arg\(32 to 63) & \$202_divisor\) & \$107_div259_arg\(64 to 95);
                      state_var1463 <= \$107_div259\;
                    end if;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("NON INT"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var1463 <= \$37_forever264958\;
                  end case;
                when pause_getII1305 =>
                  \$arr963_ptr_take\(0) := '0';
                  \$174_var\ := \$arr963_value\;
                  \$v1302\ := \$174_var\;
                  \$v1303\ := \$v1302\(0 to 3);
                  \$v1301\ := \$v1302\(4 to 67);
                  case \$v1303\ is
                  when "0001" =>
                    \$180_a\ := \$v1301\(0 to 31);
                    \$175_mult\ := \$180_a\;
                    \$108_mul260_arg\ := eclat_sub(\$108_mul260_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_mult(\$108_mul260_arg\(32 to 63) & \$175_mult\) & \$108_mul260_arg\(64 to 95);
                    state_var1463 <= \$108_mul260\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("NON INT"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var1463 <= \$37_forever264959\;
                  end case;
                when pause_getII1313 =>
                  \$arr963_ptr_take\(0) := '0';
                  \$146_var\ := \$arr963_value\;
                  \$v1310\ := \$146_var\;
                  \$v1311\ := \$v1310\(0 to 3);
                  \$v1309\ := \$v1310\(4 to 67);
                  case \$v1311\ is
                  when "0001" =>
                    \$152_a\ := \$v1309\(0 to 31);
                    \$147_sous\ := \$152_a\;
                    \$109_sub261_arg\ := eclat_sub(\$109_sub261_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_sub(\$109_sub261_arg\(32 to 63) & \$147_sous\) & \$109_sub261_arg\(64 to 95);
                    state_var1463 <= \$109_sub261\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("NON INT"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var1463 <= \$37_forever264960\;
                  end case;
                when pause_getII1321 =>
                  \$arr963_ptr_take\(0) := '0';
                  \$119_var\ := \$arr963_value\;
                  \$v1318\ := \$119_var\;
                  \$v1319\ := \$v1318\(0 to 3);
                  \$v1317\ := \$v1318\(4 to 67);
                  case \$v1319\ is
                  when "0001" =>
                    \$125_a\ := \$v1317\(0 to 31);
                    \$120_addition\ := \$125_a\;
                    \$110_add262_arg\ := eclat_sub(\$110_add262_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_add(\$110_add262_arg\(32 to 63) & \$120_addition\) & \$110_add262_arg\(64 to 95);
                    state_var1463 <= \$110_add262\;
                  when others =>
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("NON INT "));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var1463 <= \$37_forever264961\;
                  end case;
                when pause_setI1282 =>
                  \$arr962_write_request\ <= '0';
                  state_var1463 <= pause_setII1283;
                when pause_setI1326 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1327;
                when pause_setI1331 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1332;
                when pause_setI1336 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1337;
                when pause_setI1341 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1342;
                when pause_setI1346 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1347;
                when pause_setI1353 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1354;
                when pause_setI1359 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1360;
                when pause_setI1364 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1365;
                when pause_setI1369 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1370;
                when pause_setI1374 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1375;
                when pause_setI1381 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1382;
                when pause_setI1387 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1388;
                when pause_setI1392 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1393;
                when pause_setI1397 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1398;
                when pause_setI1402 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1403;
                when pause_setI1409 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1410;
                when pause_setI1414 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1415;
                when pause_setI1419 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1420;
                when pause_setI1424 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1425;
                when pause_setI1430 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1431;
                when pause_setI1435 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1436;
                when pause_setI1440 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1441;
                when pause_setI1446 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1447;
                when pause_setI1451 =>
                  \$arr965_write_request\ <= '0';
                  state_var1463 <= pause_setII1452;
                when pause_setII1283 =>
                  \$arr962_ptr_take\(0) := '0';
                  \$105_copy_args_to_heap257_arg\ := eclat_sub(\$105_copy_args_to_heap257_arg\(0 to 31) & "00000000000000000000000000000001") & \$105_copy_args_to_heap257_arg\(32 to 63) & eclat_add(\$105_copy_args_to_heap257_arg\(64 to 95) & "00000000000000000000000000000001") & \$105_copy_args_to_heap257_arg\(96 to 127) & \$105_copy_args_to_heap257_arg\(128 to 159);
                  state_var1463 <= \$105_copy_args_to_heap257\;
                when pause_setII1327 =>
                  \$arr965_ptr_take\(0) := '0';
                  result1279 := eclat_unit;
                  rdy1280 := eclat_true;
                  state_var1463 <= compute1281;
                when pause_setII1332 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1329\ := \$arr965_ptr_take\;
                  if \$v1329\(0) = '1' then
                    state_var1463 <= q_wait1328;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1325\ := eclat_unit;
                    \$arr965_ptr_write\ <= 23;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0111" & \$v1325\&"000"& X"0000000000000000";
                    state_var1463 <= pause_setI1326;
                  end if;
                when pause_setII1337 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1334\ := \$arr965_ptr_take\;
                  if \$v1334\(0) = '1' then
                    state_var1463 <= q_wait1333;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1330\ := "00000000000000000000000000000001";
                    \$arr965_ptr_write\ <= 22;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0010" & \$v1330\&X"000000000";
                    state_var1463 <= pause_setI1331;
                  end if;
                when pause_setII1342 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1339\ := \$arr965_ptr_take\;
                  if \$v1339\(0) = '1' then
                    state_var1463 <= q_wait1338;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1335\ := "00000000000000000000000000000110";
                    \$arr965_ptr_write\ <= 21;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "1010" & \$v1335\&X"000000000";
                    state_var1463 <= pause_setI1336;
                  end if;
                when pause_setII1347 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1344\ := \$arr965_ptr_take\;
                  if \$v1344\(0) = '1' then
                    state_var1463 <= q_wait1343;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1340\ := "00000000000000000000000000000000";
                    \$arr965_ptr_write\ <= 20;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0001" & \$v1340\&X"000000000";
                    state_var1463 <= pause_setI1341;
                  end if;
                when pause_setII1354 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1349\ := \$arr965_ptr_take\;
                  if \$v1349\(0) = '1' then
                    state_var1463 <= q_wait1348;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1345\ := "00000000000000000000000000000010";
                    \$arr965_ptr_write\ <= 19;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "1000" & \$v1345\&X"000000000";
                    state_var1463 <= pause_setI1346;
                  end if;
                when pause_setII1360 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1356\ := \$arr965_ptr_take\;
                  if \$v1356\(0) = '1' then
                    state_var1463 <= q_wait1355;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1350\ := eclat_unit;
                    \$v1351\ := "0001" & \$v1350\;
                    \$v1352\ := "0011" & \$v1351\&"000"& X"00000000000000";
                    \$arr965_ptr_write\ <= 18;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0101" & \$v1352\;
                    state_var1463 <= pause_setI1353;
                  end if;
                when pause_setII1365 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1362\ := \$arr965_ptr_take\;
                  if \$v1362\(0) = '1' then
                    state_var1463 <= q_wait1361;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1357\ := "00000000000000000000000000000001";
                    \$v1358\ := "0001" & \$v1357\&X"00000000";
                    \$arr965_ptr_write\ <= 17;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0101" & \$v1358\;
                    state_var1463 <= pause_setI1359;
                  end if;
                when pause_setII1370 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1367\ := \$arr965_ptr_take\;
                  if \$v1367\(0) = '1' then
                    state_var1463 <= q_wait1366;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1363\ := "00000000000000000000000000000000";
                    \$arr965_ptr_write\ <= 16;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0010" & \$v1363\&X"000000000";
                    state_var1463 <= pause_setI1364;
                  end if;
                when pause_setII1375 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1372\ := \$arr965_ptr_take\;
                  if \$v1372\(0) = '1' then
                    state_var1463 <= q_wait1371;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1368\ := X"000000" & X"16";
                    \$arr965_ptr_write\ <= 15;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "1011" & \$v1368\&X"000000000";
                    state_var1463 <= pause_setI1369;
                  end if;
                when pause_setII1382 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1377\ := \$arr965_ptr_take\;
                  if \$v1377\(0) = '1' then
                    state_var1463 <= q_wait1376;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1373\ := "00000000000000000000000000000010";
                    \$arr965_ptr_write\ <= 14;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "1000" & \$v1373\&X"000000000";
                    state_var1463 <= pause_setI1374;
                  end if;
                when pause_setII1388 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1384\ := \$arr965_ptr_take\;
                  if \$v1384\(0) = '1' then
                    state_var1463 <= q_wait1383;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1378\ := eclat_unit;
                    \$v1379\ := "0101" & \$v1378\;
                    \$v1380\ := "0011" & \$v1379\&"000"& X"00000000000000";
                    \$arr965_ptr_write\ <= 13;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0101" & \$v1380\;
                    state_var1463 <= pause_setI1381;
                  end if;
                when pause_setII1393 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1390\ := \$arr965_ptr_take\;
                  if \$v1390\(0) = '1' then
                    state_var1463 <= q_wait1389;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1385\ := "00000000000000000000000000000000";
                    \$v1386\ := "0001" & \$v1385\&X"00000000";
                    \$arr965_ptr_write\ <= 12;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0101" & \$v1386\;
                    state_var1463 <= pause_setI1387;
                  end if;
                when pause_setII1398 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1395\ := \$arr965_ptr_take\;
                  if \$v1395\(0) = '1' then
                    state_var1463 <= q_wait1394;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1391\ := "00000000000000000000000000000000";
                    \$arr965_ptr_write\ <= 11;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0010" & \$v1391\&X"000000000";
                    state_var1463 <= pause_setI1392;
                  end if;
                when pause_setII1403 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1400\ := \$arr965_ptr_take\;
                  if \$v1400\(0) = '1' then
                    state_var1463 <= q_wait1399;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1396\ := "00000000000000000000000000000001";
                    \$arr965_ptr_write\ <= 10;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0001" & \$v1396\&X"000000000";
                    state_var1463 <= pause_setI1397;
                  end if;
                when pause_setII1410 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1405\ := \$arr965_ptr_take\;
                  if \$v1405\(0) = '1' then
                    state_var1463 <= q_wait1404;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1401\ := "00000000000000000000000000000010";
                    \$arr965_ptr_write\ <= 9;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "1000" & \$v1401\&X"000000000";
                    state_var1463 <= pause_setI1402;
                  end if;
                when pause_setII1415 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1412\ := \$arr965_ptr_take\;
                  if \$v1412\(0) = '1' then
                    state_var1463 <= q_wait1411;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1406\ := eclat_unit;
                    \$v1407\ := "0000" & \$v1406\;
                    \$v1408\ := "0011" & \$v1407\&"000"& X"00000000000000";
                    \$arr965_ptr_write\ <= 8;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0101" & \$v1408\;
                    state_var1463 <= pause_setI1409;
                  end if;
                when pause_setII1420 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1417\ := \$arr965_ptr_take\;
                  if \$v1417\(0) = '1' then
                    state_var1463 <= q_wait1416;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1413\ := "00000000000000000000000000000001";
                    \$arr965_ptr_write\ <= 7;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0010" & \$v1413\&X"000000000";
                    state_var1463 <= pause_setI1414;
                  end if;
                when pause_setII1425 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1422\ := \$arr965_ptr_take\;
                  if \$v1422\(0) = '1' then
                    state_var1463 <= q_wait1421;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1418\ := "00000000000000000000000000000000";
                    \$arr965_ptr_write\ <= 6;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0010" & \$v1418\&X"000000000";
                    state_var1463 <= pause_setI1419;
                  end if;
                when pause_setII1431 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1427\ := \$arr965_ptr_take\;
                  if \$v1427\(0) = '1' then
                    state_var1463 <= q_wait1426;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1423\ := "00000000000000000000000000000001";
                    \$arr965_ptr_write\ <= 5;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0001" & \$v1423\&X"000000000";
                    state_var1463 <= pause_setI1424;
                  end if;
                when pause_setII1436 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1433\ := \$arr965_ptr_take\;
                  if \$v1433\(0) = '1' then
                    state_var1463 <= q_wait1432;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1428\ := "00000000000000000000000000000000";
                    \$v1429\ := "0001" & \$v1428\&X"00000000";
                    \$arr965_ptr_write\ <= 4;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0101" & \$v1429\;
                    state_var1463 <= pause_setI1430;
                  end if;
                when pause_setII1441 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1438\ := \$arr965_ptr_take\;
                  if \$v1438\(0) = '1' then
                    state_var1463 <= q_wait1437;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1434\ := eclat_unit;
                    \$arr965_ptr_write\ <= 3;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0000" & \$v1434\&"000"& X"0000000000000000";
                    state_var1463 <= pause_setI1435;
                  end if;
                when pause_setII1447 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1443\ := \$arr965_ptr_take\;
                  if \$v1443\(0) = '1' then
                    state_var1463 <= q_wait1442;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1439\ := "00000000000000000000000000000000";
                    \$arr965_ptr_write\ <= 2;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0001" & \$v1439\&X"000000000";
                    state_var1463 <= pause_setI1440;
                  end if;
                when pause_setII1452 =>
                  \$arr965_ptr_take\(0) := '0';
                  \$v1449\ := \$arr965_ptr_take\;
                  if \$v1449\(0) = '1' then
                    state_var1463 <= q_wait1448;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1444\ := "00000000000000000000000000001010";
                    \$v1445\ := "0001" & \$v1444\&X"00000000";
                    \$arr965_ptr_write\ <= 1;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0101" & \$v1445\;
                    state_var1463 <= pause_setI1446;
                  end if;
                when q_wait1284 =>
                  \$v1285\ := \$arr962_ptr_take\;
                  if \$v1285\(0) = '1' then
                    state_var1463 <= q_wait1284;
                  else
                    \$arr962_ptr_take\(0) := '1';
                    \$arr962_ptr_write\ <= to_integer(unsigned(\$105_copy_args_to_heap257_arg\(128 to 159)));
                    \$arr962_write_request\ <= '1';
                    \$arr962_write\ <= \$259\;
                    state_var1463 <= pause_setI1282;
                  end if;
                when q_wait1288 =>
                  \$v1289\ := \$arr963_ptr_take\;
                  if \$v1289\(0) = '1' then
                    state_var1463 <= q_wait1288;
                  else
                    \$arr963_ptr_take\(0) := '1';
                    \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$105_copy_args_to_heap257_arg\(96 to 127) & \$105_copy_args_to_heap257_arg\(0 to 31)) & "00000000000000000000000000000001")));
                    state_var1463 <= pause_getI1286;
                  end if;
                when q_wait1298 =>
                  \$v1299\ := \$arr963_ptr_take\;
                  if \$v1299\(0) = '1' then
                    state_var1463 <= q_wait1298;
                  else
                    \$arr963_ptr_take\(0) := '1';
                    \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$107_div259_arg\(64 to 95) & "00000000000000000000000000000001") & \$107_div259_arg\(0 to 31))));
                    state_var1463 <= pause_getI1296;
                  end if;
                when q_wait1306 =>
                  \$v1307\ := \$arr963_ptr_take\;
                  if \$v1307\(0) = '1' then
                    state_var1463 <= q_wait1306;
                  else
                    \$arr963_ptr_take\(0) := '1';
                    \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$108_mul260_arg\(64 to 95) & "00000000000000000000000000000001") & \$108_mul260_arg\(0 to 31))));
                    state_var1463 <= pause_getI1304;
                  end if;
                when q_wait1314 =>
                  \$v1315\ := \$arr963_ptr_take\;
                  if \$v1315\(0) = '1' then
                    state_var1463 <= q_wait1314;
                  else
                    \$arr963_ptr_take\(0) := '1';
                    \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$109_sub261_arg\(64 to 95) & "00000000000000000000000000000001") & \$109_sub261_arg\(0 to 31))));
                    state_var1463 <= pause_getI1312;
                  end if;
                when q_wait1322 =>
                  \$v1323\ := \$arr963_ptr_take\;
                  if \$v1323\(0) = '1' then
                    state_var1463 <= q_wait1322;
                  else
                    \$arr963_ptr_take\(0) := '1';
                    \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$110_add262_arg\(64 to 95) & "00000000000000000000000000000001") & \$110_add262_arg\(0 to 31))));
                    state_var1463 <= pause_getI1320;
                  end if;
                when q_wait1328 =>
                  \$v1329\ := \$arr965_ptr_take\;
                  if \$v1329\(0) = '1' then
                    state_var1463 <= q_wait1328;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1325\ := eclat_unit;
                    \$arr965_ptr_write\ <= 23;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0111" & \$v1325\&"000"& X"0000000000000000";
                    state_var1463 <= pause_setI1326;
                  end if;
                when q_wait1333 =>
                  \$v1334\ := \$arr965_ptr_take\;
                  if \$v1334\(0) = '1' then
                    state_var1463 <= q_wait1333;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1330\ := "00000000000000000000000000000001";
                    \$arr965_ptr_write\ <= 22;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0010" & \$v1330\&X"000000000";
                    state_var1463 <= pause_setI1331;
                  end if;
                when q_wait1338 =>
                  \$v1339\ := \$arr965_ptr_take\;
                  if \$v1339\(0) = '1' then
                    state_var1463 <= q_wait1338;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1335\ := "00000000000000000000000000000110";
                    \$arr965_ptr_write\ <= 21;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "1010" & \$v1335\&X"000000000";
                    state_var1463 <= pause_setI1336;
                  end if;
                when q_wait1343 =>
                  \$v1344\ := \$arr965_ptr_take\;
                  if \$v1344\(0) = '1' then
                    state_var1463 <= q_wait1343;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1340\ := "00000000000000000000000000000000";
                    \$arr965_ptr_write\ <= 20;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0001" & \$v1340\&X"000000000";
                    state_var1463 <= pause_setI1341;
                  end if;
                when q_wait1348 =>
                  \$v1349\ := \$arr965_ptr_take\;
                  if \$v1349\(0) = '1' then
                    state_var1463 <= q_wait1348;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1345\ := "00000000000000000000000000000010";
                    \$arr965_ptr_write\ <= 19;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "1000" & \$v1345\&X"000000000";
                    state_var1463 <= pause_setI1346;
                  end if;
                when q_wait1355 =>
                  \$v1356\ := \$arr965_ptr_take\;
                  if \$v1356\(0) = '1' then
                    state_var1463 <= q_wait1355;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1350\ := eclat_unit;
                    \$v1351\ := "0001" & \$v1350\;
                    \$v1352\ := "0011" & \$v1351\&"000"& X"00000000000000";
                    \$arr965_ptr_write\ <= 18;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0101" & \$v1352\;
                    state_var1463 <= pause_setI1353;
                  end if;
                when q_wait1361 =>
                  \$v1362\ := \$arr965_ptr_take\;
                  if \$v1362\(0) = '1' then
                    state_var1463 <= q_wait1361;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1357\ := "00000000000000000000000000000001";
                    \$v1358\ := "0001" & \$v1357\&X"00000000";
                    \$arr965_ptr_write\ <= 17;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0101" & \$v1358\;
                    state_var1463 <= pause_setI1359;
                  end if;
                when q_wait1366 =>
                  \$v1367\ := \$arr965_ptr_take\;
                  if \$v1367\(0) = '1' then
                    state_var1463 <= q_wait1366;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1363\ := "00000000000000000000000000000000";
                    \$arr965_ptr_write\ <= 16;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0010" & \$v1363\&X"000000000";
                    state_var1463 <= pause_setI1364;
                  end if;
                when q_wait1371 =>
                  \$v1372\ := \$arr965_ptr_take\;
                  if \$v1372\(0) = '1' then
                    state_var1463 <= q_wait1371;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1368\ := X"000000" & X"16";
                    \$arr965_ptr_write\ <= 15;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "1011" & \$v1368\&X"000000000";
                    state_var1463 <= pause_setI1369;
                  end if;
                when q_wait1376 =>
                  \$v1377\ := \$arr965_ptr_take\;
                  if \$v1377\(0) = '1' then
                    state_var1463 <= q_wait1376;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1373\ := "00000000000000000000000000000010";
                    \$arr965_ptr_write\ <= 14;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "1000" & \$v1373\&X"000000000";
                    state_var1463 <= pause_setI1374;
                  end if;
                when q_wait1383 =>
                  \$v1384\ := \$arr965_ptr_take\;
                  if \$v1384\(0) = '1' then
                    state_var1463 <= q_wait1383;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1378\ := eclat_unit;
                    \$v1379\ := "0101" & \$v1378\;
                    \$v1380\ := "0011" & \$v1379\&"000"& X"00000000000000";
                    \$arr965_ptr_write\ <= 13;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0101" & \$v1380\;
                    state_var1463 <= pause_setI1381;
                  end if;
                when q_wait1389 =>
                  \$v1390\ := \$arr965_ptr_take\;
                  if \$v1390\(0) = '1' then
                    state_var1463 <= q_wait1389;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1385\ := "00000000000000000000000000000000";
                    \$v1386\ := "0001" & \$v1385\&X"00000000";
                    \$arr965_ptr_write\ <= 12;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0101" & \$v1386\;
                    state_var1463 <= pause_setI1387;
                  end if;
                when q_wait1394 =>
                  \$v1395\ := \$arr965_ptr_take\;
                  if \$v1395\(0) = '1' then
                    state_var1463 <= q_wait1394;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1391\ := "00000000000000000000000000000000";
                    \$arr965_ptr_write\ <= 11;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0010" & \$v1391\&X"000000000";
                    state_var1463 <= pause_setI1392;
                  end if;
                when q_wait1399 =>
                  \$v1400\ := \$arr965_ptr_take\;
                  if \$v1400\(0) = '1' then
                    state_var1463 <= q_wait1399;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1396\ := "00000000000000000000000000000001";
                    \$arr965_ptr_write\ <= 10;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0001" & \$v1396\&X"000000000";
                    state_var1463 <= pause_setI1397;
                  end if;
                when q_wait1404 =>
                  \$v1405\ := \$arr965_ptr_take\;
                  if \$v1405\(0) = '1' then
                    state_var1463 <= q_wait1404;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1401\ := "00000000000000000000000000000010";
                    \$arr965_ptr_write\ <= 9;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "1000" & \$v1401\&X"000000000";
                    state_var1463 <= pause_setI1402;
                  end if;
                when q_wait1411 =>
                  \$v1412\ := \$arr965_ptr_take\;
                  if \$v1412\(0) = '1' then
                    state_var1463 <= q_wait1411;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1406\ := eclat_unit;
                    \$v1407\ := "0000" & \$v1406\;
                    \$v1408\ := "0011" & \$v1407\&"000"& X"00000000000000";
                    \$arr965_ptr_write\ <= 8;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0101" & \$v1408\;
                    state_var1463 <= pause_setI1409;
                  end if;
                when q_wait1416 =>
                  \$v1417\ := \$arr965_ptr_take\;
                  if \$v1417\(0) = '1' then
                    state_var1463 <= q_wait1416;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1413\ := "00000000000000000000000000000001";
                    \$arr965_ptr_write\ <= 7;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0010" & \$v1413\&X"000000000";
                    state_var1463 <= pause_setI1414;
                  end if;
                when q_wait1421 =>
                  \$v1422\ := \$arr965_ptr_take\;
                  if \$v1422\(0) = '1' then
                    state_var1463 <= q_wait1421;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1418\ := "00000000000000000000000000000000";
                    \$arr965_ptr_write\ <= 6;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0010" & \$v1418\&X"000000000";
                    state_var1463 <= pause_setI1419;
                  end if;
                when q_wait1426 =>
                  \$v1427\ := \$arr965_ptr_take\;
                  if \$v1427\(0) = '1' then
                    state_var1463 <= q_wait1426;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1423\ := "00000000000000000000000000000001";
                    \$arr965_ptr_write\ <= 5;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0001" & \$v1423\&X"000000000";
                    state_var1463 <= pause_setI1424;
                  end if;
                when q_wait1432 =>
                  \$v1433\ := \$arr965_ptr_take\;
                  if \$v1433\(0) = '1' then
                    state_var1463 <= q_wait1432;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1428\ := "00000000000000000000000000000000";
                    \$v1429\ := "0001" & \$v1428\&X"00000000";
                    \$arr965_ptr_write\ <= 4;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0101" & \$v1429\;
                    state_var1463 <= pause_setI1430;
                  end if;
                when q_wait1437 =>
                  \$v1438\ := \$arr965_ptr_take\;
                  if \$v1438\(0) = '1' then
                    state_var1463 <= q_wait1437;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1434\ := eclat_unit;
                    \$arr965_ptr_write\ <= 3;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0000" & \$v1434\&"000"& X"0000000000000000";
                    state_var1463 <= pause_setI1435;
                  end if;
                when q_wait1442 =>
                  \$v1443\ := \$arr965_ptr_take\;
                  if \$v1443\(0) = '1' then
                    state_var1463 <= q_wait1442;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1439\ := "00000000000000000000000000000000";
                    \$arr965_ptr_write\ <= 2;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0001" & \$v1439\&X"000000000";
                    state_var1463 <= pause_setI1440;
                  end if;
                when q_wait1448 =>
                  \$v1449\ := \$arr965_ptr_take\;
                  if \$v1449\(0) = '1' then
                    state_var1463 <= q_wait1448;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1444\ := "00000000000000000000000000001010";
                    \$v1445\ := "0001" & \$v1444\&X"00000000";
                    \$arr965_ptr_write\ <= 1;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0101" & \$v1445\;
                    state_var1463 <= pause_setI1446;
                  end if;
                when q_wait1453 =>
                  \$v1454\ := \$arr965_ptr_take\;
                  if \$v1454\(0) = '1' then
                    state_var1463 <= q_wait1453;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1450\ := eclat_unit;
                    \$arr965_ptr_write\ <= 0;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0000" & \$v1450\&"000"& X"0000000000000000";
                    state_var1463 <= pause_setI1451;
                  end if;
                when compute1281 =>
                  rdy1280 := eclat_false;
                  \$v1454\ := \$arr965_ptr_take\;
                  if \$v1454\(0) = '1' then
                    state_var1463 <= q_wait1453;
                  else
                    \$arr965_ptr_take\(0) := '1';
                    \$v1450\ := eclat_unit;
                    \$arr965_ptr_write\ <= 0;
                    \$arr965_write_request\ <= '1';
                    \$arr965_write\ <= "0000" & \$v1450\&"000"& X"0000000000000000";
                    state_var1463 <= pause_setI1451;
                  end if;
                end case;
                \$v1456\ := eclat_not(rdy1280);
                if \$v1456\(0) = '1' then
                  result1279 := eclat_unit;
                end if;
                \$v723\ := result1279 & rdy1280;
                result1276 := ""&\$v723\(1);
                rdy1277 := eclat_true;
                state_var1462 <= compute1278;
              end if;
            end case;
            \$v1459\ := eclat_not(rdy1277);
            if \$v1459\(0) = '1' then
              result1276 := eclat_false;
            end if;
            \$v722\ := result1276;
            is_loaded := result1276;
            case state_var1461 is
            when compute1273 =>
              rdy1272 := eclat_false;
              result1271 := eclat_if(is_loaded & eclat_add(\$v721\ & "00000000000000000000000000000001") & \$v721\);
              rdy1272 := eclat_true;
              state_var1461 <= compute1273;
            end case;
            \$v1275\ := eclat_not(rdy1272);
            if \$v1275\(0) = '1' then
              result1271 := "00000000000000000000000000000000";
            end if;
            \$v721\ := result1271;
            cy := result1271;
            case state_var1460 is
            when \$37_forever264932\ =>
              state_var1460 <= \$37_forever264932\;
            when \$37_forever264934\ =>
              state_var1460 <= \$87_forever264932\;
            when \$37_forever264935\ =>
              state_var1460 <= \$95_forever264932\;
            when \$37_forever264936\ =>
              state_var1460 <= \$76_forever264932\;
            when \$37_forever264937\ =>
              state_var1460 <= \$63_forever264932\;
            when \$37_forever264938\ =>
              state_var1460 <= \$37_forever264932\;
            when \$37_forever264944\ =>
              state_var1460 <= \$37_forever264932\;
            when \$37_forever264945\ =>
              state_var1460 <= \$37_forever264932\;
            when \$37_forever264946\ =>
              state_var1460 <= \$37_forever264932\;
            when \$37_forever264947\ =>
              state_var1460 <= \$37_forever264932\;
            when \$37_forever264948\ =>
              state_var1460 <= \$37_forever264932\;
            when \$37_forever264949\ =>
              state_var1460 <= \$37_forever264932\;
            when \$37_forever264950\ =>
              state_var1460 <= \$37_forever264932\;
            when \$37_forever264951\ =>
              state_var1460 <= \$37_forever264932\;
            when \$37_forever264952\ =>
              state_var1460 <= \$37_forever264932\;
            when \$37_forever264953\ =>
              state_var1460 <= \$37_forever264932\;
            when \$37_forever264954\ =>
              state_var1460 <= \$37_forever264932\;
            when \$39_copy_args_to_heap257\ =>
              \$v1025\ := eclat_eq(\$39_copy_args_to_heap257_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1025\(0) = '1' then
                \$39_copy_args_to_heap257_result\ := \$39_copy_args_to_heap257_arg\(32 to 63);
                \$v1070\ := \$arr966_ptr_take\;
                if \$v1070\(0) = '1' then
                  state_var1460 <= q_wait1069;
                else
                  \$arr966_ptr_take\(0) := '1';
                  \$arr966_ptr_write\ <= to_integer(unsigned(vm_run_code247_arg(96 to 127)));
                  \$arr966_write_request\ <= '1';
                  \$arr966_write\ <= eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127);
                  state_var1460 <= pause_setI1067;
                end if;
              else
                \$v1024\ := \$arr963_ptr_take\;
                if \$v1024\(0) = '1' then
                  state_var1460 <= q_wait1023;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$39_copy_args_to_heap257_arg\(96 to 127) & \$39_copy_args_to_heap257_arg\(0 to 31)) & "00000000000000000000000000000001")));
                  state_var1460 <= pause_getI1021;
                end if;
              end if;
            when \$40_pow258\ =>
              \$v1026\ := eclat_eq(\$40_pow258_arg\(32 to 63) & "00000000000000000000000000000000");
              if \$v1026\(0) = '1' then
                \$40_pow258_result\ := \$40_pow258_arg\(64 to 95);
                res := \$40_pow258_result\;
                \$v1125\ := \$arr963_ptr_take\;
                if \$v1125\(0) = '1' then
                  state_var1460 <= q_wait1124;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                  \$arr963_write_request\ <= '1';
                  \$arr963_write\ <= "0001" & res&X"00000000";
                  state_var1460 <= pause_setI1122;
                end if;
              else
                \$40_pow258_arg\ := \$40_pow258_arg\(0 to 31) & eclat_sub(\$40_pow258_arg\(32 to 63) & "00000000000000000000000000000001") & eclat_mult(\$40_pow258_arg\(64 to 95) & \$40_pow258_arg\(0 to 31));
                state_var1460 <= \$40_pow258\;
              end if;
            when \$41_div259\ =>
              \$v1035\ := eclat_eq(\$41_div259_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1035\(0) = '1' then
                \$41_div259_result\ := \$41_div259_arg\(32 to 63);
                res := \$41_div259_result\;
                \$v1144\ := \$arr963_ptr_take\;
                if \$v1144\(0) = '1' then
                  state_var1460 <= q_wait1143;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                  \$arr963_write_request\ <= '1';
                  \$arr963_write\ <= "0001" & res&X"00000000";
                  state_var1460 <= pause_setI1141;
                end if;
              else
                \$v1034\ := \$arr963_ptr_take\;
                if \$v1034\(0) = '1' then
                  state_var1460 <= q_wait1033;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$41_div259_arg\(64 to 95) & "00000000000000000000000000000001") & \$41_div259_arg\(0 to 31))));
                  state_var1460 <= pause_getI1031;
                end if;
              end if;
            when \$42_mul260\ =>
              \$v1043\ := eclat_eq(\$42_mul260_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1043\(0) = '1' then
                \$42_mul260_result\ := \$42_mul260_arg\(32 to 63);
                res := \$42_mul260_result\;
                \$v1156\ := \$arr963_ptr_take\;
                if \$v1156\(0) = '1' then
                  state_var1460 <= q_wait1155;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                  \$arr963_write_request\ <= '1';
                  \$arr963_write\ <= "0001" & res&X"00000000";
                  state_var1460 <= pause_setI1153;
                end if;
              else
                \$v1042\ := \$arr963_ptr_take\;
                if \$v1042\(0) = '1' then
                  state_var1460 <= q_wait1041;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$42_mul260_arg\(64 to 95) & "00000000000000000000000000000001") & \$42_mul260_arg\(0 to 31))));
                  state_var1460 <= pause_getI1039;
                end if;
              end if;
            when \$43_sub261\ =>
              \$v1051\ := eclat_eq(\$43_sub261_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1051\(0) = '1' then
                \$43_sub261_result\ := \$43_sub261_arg\(32 to 63);
                resultat := \$43_sub261_result\;
                \$v1161\ := \$arr963_ptr_take\;
                if \$v1161\(0) = '1' then
                  state_var1460 <= q_wait1160;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$v1157\ := eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat);
                  \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                  \$arr963_write_request\ <= '1';
                  \$arr963_write\ <= "0001" & \$v1157\&X"00000000";
                  state_var1460 <= pause_setI1158;
                end if;
              else
                \$v1050\ := \$arr963_ptr_take\;
                if \$v1050\(0) = '1' then
                  state_var1460 <= q_wait1049;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$43_sub261_arg\(64 to 95) & "00000000000000000000000000000001") & \$43_sub261_arg\(0 to 31))));
                  state_var1460 <= pause_getI1047;
                end if;
              end if;
            when \$44_add262\ =>
              \$v1059\ := eclat_eq(\$44_add262_arg\(0 to 31) & "00000000000000000000000000000000");
              if \$v1059\(0) = '1' then
                \$44_add262_result\ := \$44_add262_arg\(32 to 63);
                res := \$44_add262_result\;
                \$v1173\ := \$arr963_ptr_take\;
                if \$v1173\(0) = '1' then
                  state_var1460 <= q_wait1172;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                  \$arr963_write_request\ <= '1';
                  \$arr963_write\ <= "0001" & res&X"00000000";
                  state_var1460 <= pause_setI1170;
                end if;
              else
                \$v1058\ := \$arr963_ptr_take\;
                if \$v1058\(0) = '1' then
                  state_var1460 <= q_wait1057;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$44_add262_arg\(64 to 95) & "00000000000000000000000000000001") & \$44_add262_arg\(0 to 31))));
                  state_var1460 <= pause_getI1055;
                end if;
              end if;
            when \$63_forever264932\ =>
              state_var1460 <= \$63_forever264932\;
            when \$76_forever264932\ =>
              state_var1460 <= \$76_forever264932\;
            when \$87_forever264932\ =>
              state_var1460 <= \$87_forever264932\;
            when \$95_forever264932\ =>
              state_var1460 <= \$95_forever264932\;
            when forever263933 =>
              state_var1460 <= forever263933;
            when forever263939 =>
              state_var1460 <= forever263933;
            when forever263940 =>
              state_var1460 <= forever263933;
            when forever263941 =>
              state_var1460 <= forever263933;
            when forever263942 =>
              state_var1460 <= forever263933;
            when forever263943 =>
              state_var1460 <= forever263933;
            when pause_getI1021 =>
              state_var1460 <= pause_getII1022;
            when pause_getI1031 =>
              state_var1460 <= pause_getII1032;
            when pause_getI1039 =>
              state_var1460 <= pause_getII1040;
            when pause_getI1047 =>
              state_var1460 <= pause_getII1048;
            when pause_getI1055 =>
              state_var1460 <= pause_getII1056;
            when pause_getI1093 =>
              state_var1460 <= pause_getII1094;
            when pause_getI1097 =>
              state_var1460 <= pause_getII1098;
            when pause_getI1110 =>
              state_var1460 <= pause_getII1111;
            when pause_getI1117 =>
              state_var1460 <= pause_getII1118;
            when pause_getI1129 =>
              state_var1460 <= pause_getII1130;
            when pause_getI1136 =>
              state_var1460 <= pause_getII1137;
            when pause_getI1148 =>
              state_var1460 <= pause_getII1149;
            when pause_getI1165 =>
              state_var1460 <= pause_getII1166;
            when pause_getI1178 =>
              state_var1460 <= pause_getII1179;
            when pause_getI1185 =>
              state_var1460 <= pause_getII1186;
            when pause_getI1192 =>
              state_var1460 <= pause_getII1193;
            when pause_getI1200 =>
              state_var1460 <= pause_getII1201;
            when pause_getI1213 =>
              state_var1460 <= pause_getII1214;
            when pause_getI1217 =>
              state_var1460 <= pause_getII1218;
            when pause_getI1225 =>
              state_var1460 <= pause_getII1226;
            when pause_getI1236 =>
              state_var1460 <= pause_getII1237;
            when pause_getI1249 =>
              state_var1460 <= pause_getII1250;
            when pause_getI1257 =>
              state_var1460 <= pause_getII1258;
            when pause_getI1263 =>
              state_var1460 <= pause_getII1264;
            when pause_getII1022 =>
              \$arr963_ptr_take\(0) := '0';
              \$v13\ := \$arr963_value\;
              \$v1020\ := \$arr962_ptr_take\;
              if \$v1020\(0) = '1' then
                state_var1460 <= q_wait1019;
              else
                \$arr962_ptr_take\(0) := '1';
                \$arr962_ptr_write\ <= to_integer(unsigned(\$39_copy_args_to_heap257_arg\(128 to 159)));
                \$arr962_write_request\ <= '1';
                \$arr962_write\ <= \$v13\;
                state_var1460 <= pause_setI1017;
              end if;
            when pause_getII1032 =>
              \$arr963_ptr_take\(0) := '0';
              \$v70\ := \$arr963_value\;
              \$v1029\ := \$v70\;
              \$v1030\ := \$v1029\(0 to 3);
              \$v1028\ := \$v1029\(4 to 67);
              case \$v1030\ is
              when "0001" =>
                \$91_a\ := \$v1028\(0 to 31);
                divisor := \$91_a\;
                \$v1027\ := eclat_eq(divisor & "00000000000000000000000000000000");
                if \$v1027\(0) = '1' then
                  eclat_print_string(of_string("fatal error: "));
                  
                  eclat_print_string(of_string("Div par zero impossible"));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var1460 <= \$37_forever264934\;
                else
                  \$41_div259_arg\ := eclat_sub(\$41_div259_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_div(\$41_div259_arg\(32 to 63) & divisor) & \$41_div259_arg\(64 to 95);
                  state_var1460 <= \$41_div259\;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("NON INT"));
                
                eclat_print_newline(eclat_unit);
                
                state_var1460 <= \$37_forever264935\;
              end case;
            when pause_getII1040 =>
              \$arr963_ptr_take\(0) := '0';
              \$71_var\ := \$arr963_value\;
              \$v1037\ := \$71_var\;
              \$v1038\ := \$v1037\(0 to 3);
              \$v1036\ := \$v1037\(4 to 67);
              case \$v1038\ is
              when "0001" =>
                \$72_a\ := \$v1036\(0 to 31);
                mult := \$72_a\;
                \$42_mul260_arg\ := eclat_sub(\$42_mul260_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_mult(\$42_mul260_arg\(32 to 63) & mult) & \$42_mul260_arg\(64 to 95);
                state_var1460 <= \$42_mul260\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("NON INT"));
                
                eclat_print_newline(eclat_unit);
                
                state_var1460 <= \$37_forever264936\;
              end case;
            when pause_getII1048 =>
              \$arr963_ptr_take\(0) := '0';
              \$58_var\ := \$arr963_value\;
              \$v1045\ := \$58_var\;
              \$v1046\ := \$v1045\(0 to 3);
              \$v1044\ := \$v1045\(4 to 67);
              case \$v1046\ is
              when "0001" =>
                \$59_a\ := \$v1044\(0 to 31);
                sous := \$59_a\;
                \$43_sub261_arg\ := eclat_sub(\$43_sub261_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_sub(\$43_sub261_arg\(32 to 63) & sous) & \$43_sub261_arg\(64 to 95);
                state_var1460 <= \$43_sub261\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("NON INT"));
                
                eclat_print_newline(eclat_unit);
                
                state_var1460 <= \$37_forever264937\;
              end case;
            when pause_getII1056 =>
              \$arr963_ptr_take\(0) := '0';
              var := \$arr963_value\;
              \$v1053\ := var;
              \$v1054\ := \$v1053\(0 to 3);
              \$v1052\ := \$v1053\(4 to 67);
              case \$v1054\ is
              when "0001" =>
                a := \$v1052\(0 to 31);
                addition := a;
                \$44_add262_arg\ := eclat_sub(\$44_add262_arg\(0 to 31) & "00000000000000000000000000000001") & eclat_add(\$44_add262_arg\(32 to 63) & addition) & \$44_add262_arg\(64 to 95);
                state_var1460 <= \$44_add262\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("NON INT "));
                
                eclat_print_newline(eclat_unit);
                
                state_var1460 <= \$37_forever264938\;
              end case;
            when pause_getII1094 =>
              \$arr963_ptr_take\(0) := '0';
              e2 := \$arr963_value\;
              \$v1091\ := e1;
              \$v1092\ := \$v1091\(0 to 3);
              \$v1081\ := \$v1091\(4 to 67);
              case \$v1092\ is
              when "0010" =>
                \$v1083\ := e2;
                \$v1084\ := \$v1083\(0 to 3);
                \$v1082\ := \$v1083\(4 to 67);
                case \$v1084\ is
                when "0010" =>
                  verif := eclat_true;
                  \$v1080\ := \$arr963_ptr_take\;
                  if \$v1080\(0) = '1' then
                    state_var1460 <= q_wait1079;
                  else
                    \$arr963_ptr_take\(0) := '1';
                    \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & n)));
                    \$arr963_write_request\ <= '1';
                    \$arr963_write\ <= "0000" & verif&"000"& X"000000000000000";
                    state_var1460 <= pause_setI1077;
                  end if;
                when others =>
                  eclat_print_string(of_string("Pas pareil\n"));
                  
                  eclat_print_string(of_string("(exit) bye bye."));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var1460 <= forever263941;
                end case;
              when "0000" =>
                a1 := \$v1081\(0 to 0);
                \$v1086\ := e2;
                \$v1087\ := \$v1086\(0 to 3);
                \$v1085\ := \$v1086\(4 to 67);
                case \$v1087\ is
                when "0000" =>
                  b2 := \$v1085\(0 to 0);
                  verif := eclat_if(a1 & eclat_if(b2 & eclat_true & eclat_false) & 
                           eclat_if(b2 & eclat_false & eclat_true));
                  \$v1080\ := \$arr963_ptr_take\;
                  if \$v1080\(0) = '1' then
                    state_var1460 <= q_wait1079;
                  else
                    \$arr963_ptr_take\(0) := '1';
                    \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & n)));
                    \$arr963_write_request\ <= '1';
                    \$arr963_write\ <= "0000" & verif&"000"& X"000000000000000";
                    state_var1460 <= pause_setI1077;
                  end if;
                when others =>
                  eclat_print_string(of_string("Les 2 sont pas BOOL\n"));
                  
                  eclat_print_string(of_string("(exit) bye bye."));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var1460 <= forever263942;
                end case;
              when "0001" =>
                a := \$v1081\(0 to 31);
                \$v1089\ := e2;
                \$v1090\ := \$v1089\(0 to 3);
                \$v1088\ := \$v1089\(4 to 67);
                case \$v1090\ is
                when "0001" =>
                  b := \$v1088\(0 to 31);
                  verif := eclat_eq(a & b);
                  \$v1080\ := \$arr963_ptr_take\;
                  if \$v1080\(0) = '1' then
                    state_var1460 <= q_wait1079;
                  else
                    \$arr963_ptr_take\(0) := '1';
                    \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & n)));
                    \$arr963_write_request\ <= '1';
                    \$arr963_write\ <= "0000" & verif&"000"& X"000000000000000";
                    state_var1460 <= pause_setI1077;
                  end if;
                when others =>
                  eclat_print_string(of_string("Les 2 sont pas INT\n"));
                  
                  eclat_print_string(of_string("(exit) bye bye."));
                  
                  eclat_print_newline(eclat_unit);
                  
                  state_var1460 <= forever263943;
                end case;
              when others =>
                eclat_print_string(of_string("Erreur \n"));
                
                eclat_print_string(of_string("(exit) bye bye."));
                
                eclat_print_newline(eclat_unit);
                
                state_var1460 <= forever263940;
              end case;
            when pause_getII1098 =>
              \$arr963_ptr_take\(0) := '0';
              e1 := \$arr963_value\;
              \$v1096\ := \$arr963_ptr_take\;
              if \$v1096\(0) = '1' then
                state_var1460 <= q_wait1095;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000011")));
                state_var1460 <= pause_getI1093;
              end if;
            when pause_getII1111 =>
              \$arr963_ptr_take\(0) := '0';
              \$v43\ := \$arr963_value\;
              \$v1108\ := \$v43\;
              \$v1109\ := \$v1108\(0 to 3);
              \$v1107\ := \$v1108\(4 to 67);
              case \$v1109\ is
              when "0001" =>
                a := \$v1107\(0 to 31);
                b := a;
                \$v1106\ := \$arr963_ptr_take\;
                if \$v1106\(0) = '1' then
                  state_var1460 <= q_wait1105;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$v1102\ := eclat_gt(a & b);
                  \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                  \$arr963_write_request\ <= '1';
                  \$arr963_write\ <= "0000" & \$v1102\&"000"& X"000000000000000";
                  state_var1460 <= pause_setI1103;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("NON INT"));
                
                eclat_print_newline(eclat_unit);
                
                state_var1460 <= \$37_forever264945\;
              end case;
            when pause_getII1118 =>
              \$arr963_ptr_take\(0) := '0';
              \$v41\ := \$arr963_value\;
              \$v1115\ := \$v41\;
              \$v1116\ := \$v1115\(0 to 3);
              \$v1114\ := \$v1115\(4 to 67);
              case \$v1116\ is
              when "0001" =>
                a := \$v1114\(0 to 31);
                a := a;
                \$v1113\ := \$arr963_ptr_take\;
                if \$v1113\(0) = '1' then
                  state_var1460 <= q_wait1112;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000010")));
                  state_var1460 <= pause_getI1110;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("NON INT"));
                
                eclat_print_newline(eclat_unit);
                
                state_var1460 <= \$37_forever264946\;
              end case;
            when pause_getII1130 =>
              \$arr963_ptr_take\(0) := '0';
              \$v54\ := \$arr963_value\;
              \$v1127\ := \$v54\;
              \$v1128\ := \$v1127\(0 to 3);
              \$v1126\ := \$v1127\(4 to 67);
              case \$v1128\ is
              when "0001" =>
                a := \$v1126\(0 to 31);
                puissance := a;
                \$40_pow258_arg\ := i & puissance & "00000000000000000000000000000001";
                state_var1460 <= \$40_pow258\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("NON INT"));
                
                eclat_print_newline(eclat_unit);
                
                state_var1460 <= \$37_forever264948\;
              end case;
            when pause_getII1137 =>
              \$arr963_ptr_take\(0) := '0';
              \$v52\ := \$arr963_value\;
              \$v1134\ := \$v52\;
              \$v1135\ := \$v1134\(0 to 3);
              \$v1133\ := \$v1134\(4 to 67);
              case \$v1135\ is
              when "0001" =>
                a := \$v1133\(0 to 31);
                i := a;
                \$v1132\ := \$arr963_ptr_take\;
                if \$v1132\(0) = '1' then
                  state_var1460 <= q_wait1131;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000010")));
                  state_var1460 <= pause_getI1129;
                end if;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("NON INT"));
                
                eclat_print_newline(eclat_unit);
                
                state_var1460 <= \$37_forever264949\;
              end case;
            when pause_getII1149 =>
              \$arr963_ptr_take\(0) := '0';
              \$v78\ := \$arr963_value\;
              \$v1146\ := \$v78\;
              \$v1147\ := \$v1146\(0 to 3);
              \$v1145\ := \$v1146\(4 to 67);
              case \$v1147\ is
              when "0001" =>
                a := \$v1145\(0 to 31);
                valeur_depart := a;
                \$41_div259_arg\ := eclat_sub(n & "00000000000000000000000000000001") & valeur_depart & vm_run_code247_arg(0 to 31);
                state_var1460 <= \$41_div259\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("NON INT"));
                
                eclat_print_newline(eclat_unit);
                
                state_var1460 <= \$37_forever264951\;
              end case;
            when pause_getII1166 =>
              \$arr963_ptr_take\(0) := '0';
              \$v111\ := \$arr963_value\;
              \$v1163\ := \$v111\;
              \$v1164\ := \$v1163\(0 to 3);
              \$v1162\ := \$v1163\(4 to 67);
              case \$v1164\ is
              when "0001" =>
                a := \$v1162\(0 to 31);
                valeur_depart := a;
                \$43_sub261_arg\ := eclat_sub(n & "00000000000000000000000000000001") & valeur_depart & vm_run_code247_arg(0 to 31);
                state_var1460 <= \$43_sub261\;
              when others =>
                eclat_print_string(of_string("fatal error: "));
                
                eclat_print_string(of_string("NON INT"));
                
                eclat_print_newline(eclat_unit);
                
                state_var1460 <= \$37_forever264953\;
              end case;
            when pause_getII1179 =>
              \$arr963_ptr_take\(0) := '0';
              \value\ := \$arr963_value\;
              \$v1176\ := \value\;
              \$v1177\ := \$v1176\(0 to 3);
              \$v1062\ := \$v1176\(4 to 67);
              case \$v1177\ is
              when "0100" =>
                \$v760\ := \$v1062\(0 to 63);
                \$v1075\ := \$arr962_ptr_take\;
                if \$v1075\(0) = '1' then
                  state_var1460 <= q_wait1074;
                else
                  \$arr962_ptr_take\(0) := '1';
                  \$v1071\ := vm_run_code247_arg(32 to 63);
                  \$arr962_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_add(eclat_add(vm_run_code247_arg(160 to 191) & n) & "00000000000000000000000000000001") & "00000000000000000000000000000001")));
                  \$arr962_write_request\ <= '1';
                  \$arr962_write\ <= "0001" & \$v1071\&X"00000000";
                  state_var1460 <= pause_setI1072;
                end if;
              when "0011" =>
                p := \$v1062\(0 to 4);
                \$v1174\ := p;
                \$v1175\ := \$v1174\(0 to 3);
                \$v1076\ := ""&\$v1174\(4);
                case \$v1175\ is
                when "0101" =>
                  \$v1101\ := eclat_neq(n & "00000000000000000000000000000010");
                  if \$v1101\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("Exact 2 args"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var1460 <= \$37_forever264944\;
                  else
                    \$v1100\ := \$arr963_ptr_take\;
                    if \$v1100\(0) = '1' then
                      state_var1460 <= q_wait1099;
                    else
                      \$arr963_ptr_take\(0) := '1';
                      \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000010")));
                      state_var1460 <= pause_getI1097;
                    end if;
                  end if;
                when "0110" =>
                  \$v1121\ := eclat_neq(n & "00000000000000000000000000000010");
                  if \$v1121\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("Exact 2 args"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var1460 <= \$37_forever264947\;
                  else
                    \$v1120\ := \$arr963_ptr_take\;
                    if \$v1120\(0) = '1' then
                      state_var1460 <= q_wait1119;
                    else
                      \$arr963_ptr_take\(0) := '1';
                      \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000011")));
                      state_var1460 <= pause_getI1117;
                    end if;
                  end if;
                when "0100" =>
                  \$v1140\ := eclat_neq(n & "00000000000000000000000000000010");
                  if \$v1140\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("Exact 2 args"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var1460 <= \$37_forever264950\;
                  else
                    \$v1139\ := \$arr963_ptr_take\;
                    if \$v1139\(0) = '1' then
                      state_var1460 <= q_wait1138;
                    else
                      \$arr963_ptr_take\(0) := '1';
                      \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000011")));
                      state_var1460 <= pause_getI1136;
                    end if;
                  end if;
                when "0011" =>
                  \$v1152\ := eclat_lt(n & "00000000000000000000000000000001");
                  if \$v1152\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("Min 2 args"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var1460 <= \$37_forever264952\;
                  else
                    \$v1151\ := \$arr963_ptr_take\;
                    if \$v1151\(0) = '1' then
                      state_var1460 <= q_wait1150;
                    else
                      \$arr963_ptr_take\(0) := '1';
                      \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                      state_var1460 <= pause_getI1148;
                    end if;
                  end if;
                when "0010" =>
                  \$42_mul260_arg\ := n & "00000000000000000000000000000001" & vm_run_code247_arg(0 to 31);
                  state_var1460 <= \$42_mul260\;
                when "0001" =>
                  \$v1169\ := eclat_lt(n & "00000000000000000000000000000010");
                  if \$v1169\(0) = '1' then
                    eclat_print_string(of_string("fatal error: "));
                    
                    eclat_print_string(of_string("Min 2 args"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    state_var1460 <= \$37_forever264954\;
                  else
                    \$v1168\ := \$arr963_ptr_take\;
                    if \$v1168\(0) = '1' then
                      state_var1460 <= q_wait1167;
                    else
                      \$arr963_ptr_take\(0) := '1';
                      \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                      state_var1460 <= pause_getI1165;
                    end if;
                  end if;
                when "0000" =>
                  \$44_add262_arg\ := n & "00000000000000000000000000000000" & vm_run_code247_arg(0 to 31);
                  state_var1460 <= \$44_add262\;
                when others =>
                  \$v752\ := vm_run_code247_arg(0 to 293);
                  \$v1060\ := ""&\$v752\(293);
                  if \$v1060\(0) = '1' then
                    vm_run_code247_result := eclat_unit;
                    result1014 := vm_run_code247_result;
                    rdy1015 := eclat_true;
                    state_var1460 <= compute1016;
                  else
                    vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                    state_var1460 <= vm_run_code247;
                  end if;
                end case;
              when others =>
                \$v752\ := vm_run_code247_arg(0 to 293);
                \$v1060\ := ""&\$v752\(293);
                if \$v1060\(0) = '1' then
                  vm_run_code247_result := eclat_unit;
                  result1014 := vm_run_code247_result;
                  rdy1015 := eclat_true;
                  state_var1460 <= compute1016;
                else
                  vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                  state_var1460 <= vm_run_code247;
                end if;
              end case;
            when pause_getII1186 =>
              \$arr963_ptr_take\(0) := '0';
              var := \$arr963_value\;
              \$v1183\ := var;
              \$v1184\ := \$v1183\(0 to 3);
              \$v1182\ := \$v1183\(4 to 67);
              case \$v1184\ is
              when "0000" =>
                x := \$v1182\(0 to 0);
                jfalse := x;
                \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & 
                eclat_if(jfalse & vm_run_code247_arg(64 to 95) & eclat_sub(l & "00000000000000000000000000000001")) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
                \$v1060\ := ""&\$v752\(293);
                if \$v1060\(0) = '1' then
                  vm_run_code247_result := eclat_unit;
                  result1014 := vm_run_code247_result;
                  rdy1015 := eclat_true;
                  state_var1460 <= compute1016;
                else
                  vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                  state_var1460 <= vm_run_code247;
                end if;
              when others =>
                jfalse := eclat_false;
                \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & 
                eclat_if(jfalse & vm_run_code247_arg(64 to 95) & eclat_sub(l & "00000000000000000000000000000001")) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
                \$v1060\ := ""&\$v752\(293);
                if \$v1060\(0) = '1' then
                  vm_run_code247_result := eclat_unit;
                  result1014 := vm_run_code247_result;
                  rdy1015 := eclat_true;
                  state_var1460 <= compute1016;
                else
                  vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                  state_var1460 <= vm_run_code247;
                end if;
              end case;
            when pause_getII1193 =>
              \$arr963_ptr_take\(0) := '0';
              var := \$arr963_value\;
              \$v1190\ := var;
              \$v1191\ := \$v1190\(0 to 3);
              \$v1189\ := \$v1190\(4 to 67);
              case \$v1191\ is
              when "0000" =>
                x := \$v1189\(0 to 0);
                jtrue := x;
                \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & 
                eclat_if(jtrue & eclat_sub(\$17_l\ & "00000000000000000000000000000001") & vm_run_code247_arg(64 to 95)) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
                \$v1060\ := ""&\$v752\(293);
                if \$v1060\(0) = '1' then
                  vm_run_code247_result := eclat_unit;
                  result1014 := vm_run_code247_result;
                  rdy1015 := eclat_true;
                  state_var1460 <= compute1016;
                else
                  vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                  state_var1460 <= vm_run_code247;
                end if;
              when others =>
                jtrue := eclat_false;
                \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & 
                eclat_if(jtrue & eclat_sub(\$17_l\ & "00000000000000000000000000000001") & vm_run_code247_arg(64 to 95)) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
                \$v1060\ := ""&\$v752\(293);
                if \$v1060\(0) = '1' then
                  vm_run_code247_result := eclat_unit;
                  result1014 := vm_run_code247_result;
                  rdy1015 := eclat_true;
                  state_var1460 <= compute1016;
                else
                  vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                  state_var1460 <= vm_run_code247;
                end if;
              end case;
            when pause_getII1201 =>
              \$arr963_ptr_take\(0) := '0';
              var := \$arr963_value\;
              \$v1199\ := \$arr962_ptr_take\;
              if \$v1199\(0) = '1' then
                state_var1460 <= q_wait1198;
              else
                \$arr962_ptr_take\(0) := '1';
                \$arr962_ptr_write\ <= to_integer(unsigned(eclat_add(vm_run_code247_arg(32 to 63) & i)));
                \$arr962_write_request\ <= '1';
                \$arr962_write\ <= var;
                state_var1460 <= pause_setI1196;
              end if;
            when pause_getII1214 =>
              \$arr963_ptr_take\(0) := '0';
              \$v151\ := \$arr963_value\;
              \$v1212\ := \$arr963_ptr_take\;
              if \$v1212\(0) = '1' then
                state_var1460 <= q_wait1211;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr_write\ <= to_integer(unsigned(\$v843\(0 to 31)));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= \$v151\;
                state_var1460 <= pause_setI1209;
              end if;
            when pause_getII1218 =>
              \$arr966_ptr_take\(0) := '0';
              \$v843\ := \$arr966_value\;
              \$v1216\ := \$arr963_ptr_take\;
              if \$v1216\(0) = '1' then
                state_var1460 <= q_wait1215;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001")));
                state_var1460 <= pause_getI1213;
              end if;
            when pause_getII1226 =>
              \$arr962_ptr_take\(0) := '0';
              temp := \$arr962_value\;
              \$v1224\ := \$arr963_ptr_take\;
              if \$v1224\(0) = '1' then
                state_var1460 <= q_wait1223;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr_write\ <= to_integer(unsigned(vm_run_code247_arg(0 to 31)));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= temp;
                state_var1460 <= pause_setI1221;
              end if;
            when pause_getII1237 =>
              \$arr963_ptr_take\(0) := '0';
              \$v165\ := \$arr963_value\;
              \$v1234\ := \$v165\;
              \$v1235\ := \$v1234\(0 to 3);
              \$v1229\ := \$v1234\(4 to 67);
              case \$v1235\ is
              when "0100" =>
                eclat_print_string(of_string("fermeture"));
                
                \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & eclat_true;
                \$v1060\ := ""&\$v752\(293);
                if \$v1060\(0) = '1' then
                  vm_run_code247_result := eclat_unit;
                  result1014 := vm_run_code247_result;
                  rdy1015 := eclat_true;
                  state_var1460 <= compute1016;
                else
                  vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                  state_var1460 <= vm_run_code247;
                end if;
              when "0011" =>
                p := \$v1229\(0 to 4);
                \$v1231\ := p;
                \$v1232\ := \$v1231\(0 to 3);
                \$v1230\ := ""&\$v1231\(4);
                case \$v1232\ is
                when "0110" =>
                  eclat_print_string(of_string("<"));
                  
                  \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & eclat_true;
                  \$v1060\ := ""&\$v752\(293);
                  if \$v1060\(0) = '1' then
                    vm_run_code247_result := eclat_unit;
                    result1014 := vm_run_code247_result;
                    rdy1015 := eclat_true;
                    state_var1460 <= compute1016;
                  else
                    vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                    state_var1460 <= vm_run_code247;
                  end if;
                when "0101" =>
                  eclat_print_string(of_string("=="));
                  
                  \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & eclat_true;
                  \$v1060\ := ""&\$v752\(293);
                  if \$v1060\(0) = '1' then
                    vm_run_code247_result := eclat_unit;
                    result1014 := vm_run_code247_result;
                    rdy1015 := eclat_true;
                    state_var1460 <= compute1016;
                  else
                    vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                    state_var1460 <= vm_run_code247;
                  end if;
                when "0100" =>
                  eclat_print_string(of_string("pow"));
                  
                  \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & eclat_true;
                  \$v1060\ := ""&\$v752\(293);
                  if \$v1060\(0) = '1' then
                    vm_run_code247_result := eclat_unit;
                    result1014 := vm_run_code247_result;
                    rdy1015 := eclat_true;
                    state_var1460 <= compute1016;
                  else
                    vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                    state_var1460 <= vm_run_code247;
                  end if;
                when "0011" =>
                  eclat_print_string(of_string("/"));
                  
                  \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & eclat_true;
                  \$v1060\ := ""&\$v752\(293);
                  if \$v1060\(0) = '1' then
                    vm_run_code247_result := eclat_unit;
                    result1014 := vm_run_code247_result;
                    rdy1015 := eclat_true;
                    state_var1460 <= compute1016;
                  else
                    vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                    state_var1460 <= vm_run_code247;
                  end if;
                when "0010" =>
                  eclat_print_string(of_string("*"));
                  
                  \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & eclat_true;
                  \$v1060\ := ""&\$v752\(293);
                  if \$v1060\(0) = '1' then
                    vm_run_code247_result := eclat_unit;
                    result1014 := vm_run_code247_result;
                    rdy1015 := eclat_true;
                    state_var1460 <= compute1016;
                  else
                    vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                    state_var1460 <= vm_run_code247;
                  end if;
                when "0001" =>
                  eclat_print_string(of_string("-"));
                  
                  \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & eclat_true;
                  \$v1060\ := ""&\$v752\(293);
                  if \$v1060\(0) = '1' then
                    vm_run_code247_result := eclat_unit;
                    result1014 := vm_run_code247_result;
                    rdy1015 := eclat_true;
                    state_var1460 <= compute1016;
                  else
                    vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                    state_var1460 <= vm_run_code247;
                  end if;
                when "0000" =>
                  eclat_print_string(of_string("+"));
                  
                  \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & eclat_true;
                  \$v1060\ := ""&\$v752\(293);
                  if \$v1060\(0) = '1' then
                    vm_run_code247_result := eclat_unit;
                    result1014 := vm_run_code247_result;
                    rdy1015 := eclat_true;
                    state_var1460 <= compute1016;
                  else
                    vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                    state_var1460 <= vm_run_code247;
                  end if;
                when others =>
                  
                end case;
              when "0010" =>
                eclat_print_string(of_string("nil"));
                
                \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & eclat_true;
                \$v1060\ := ""&\$v752\(293);
                if \$v1060\(0) = '1' then
                  vm_run_code247_result := eclat_unit;
                  result1014 := vm_run_code247_result;
                  rdy1015 := eclat_true;
                  state_var1460 <= compute1016;
                else
                  vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                  state_var1460 <= vm_run_code247;
                end if;
              when "0001" =>
                \$33_n\ := \$v1229\(0 to 31);
                eclat_print_int(\$33_n\);
                
                \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & eclat_true;
                \$v1060\ := ""&\$v752\(293);
                if \$v1060\(0) = '1' then
                  vm_run_code247_result := eclat_unit;
                  result1014 := vm_run_code247_result;
                  rdy1015 := eclat_true;
                  state_var1460 <= compute1016;
                else
                  vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                  state_var1460 <= vm_run_code247;
                end if;
              when "0000" =>
                \$34_b\ := \$v1229\(0 to 0);
                \$v1233\ := \$34_b\;
                if \$v1233\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & eclat_true;
                  \$v1060\ := ""&\$v752\(293);
                  if \$v1060\(0) = '1' then
                    vm_run_code247_result := eclat_unit;
                    result1014 := vm_run_code247_result;
                    rdy1015 := eclat_true;
                    state_var1460 <= compute1016;
                  else
                    vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                    state_var1460 <= vm_run_code247;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & eclat_true;
                  \$v1060\ := ""&\$v752\(293);
                  if \$v1060\(0) = '1' then
                    vm_run_code247_result := eclat_unit;
                    result1014 := vm_run_code247_result;
                    rdy1015 := eclat_true;
                    state_var1460 <= compute1016;
                  else
                    vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                    state_var1460 <= vm_run_code247;
                  end if;
                end if;
              when others =>
                
              end case;
            when pause_getII1250 =>
              \$arr964_ptr_take\(0) := '0';
              \$v170\ := \$arr964_value\;
              \$v1248\ := \$arr963_ptr_take\;
              if \$v1248\(0) = '1' then
                state_var1460 <= q_wait1247;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr_write\ <= to_integer(unsigned(vm_run_code247_arg(0 to 31)));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= \$v170\;
                state_var1460 <= pause_setI1245;
              end if;
            when pause_getII1258 =>
              \$arr963_ptr_take\(0) := '0';
              \$v174\ := \$arr963_value\;
              \$v1256\ := \$arr964_ptr_take\;
              if \$v1256\(0) = '1' then
                state_var1460 <= q_wait1255;
              else
                \$arr964_ptr_take\(0) := '1';
                \$arr964_ptr_write\ <= to_integer(unsigned(\$22_i\));
                \$arr964_write_request\ <= '1';
                \$arr964_write\ <= \$v174\;
                state_var1460 <= pause_setI1253;
              end if;
            when pause_getII1264 =>
              \$arr965_ptr_take\(0) := '0';
              instr := \$arr965_value\;
              \$v1261\ := instr;
              \$v1262\ := \$v1261\(0 to 3);
              \$v1061\ := \$v1261\(4 to 71);
              case \$v1262\ is
              when "1000" =>
                n := \$v1061\(0 to 31);
                \$v1181\ := \$arr963_ptr_take\;
                if \$v1181\(0) = '1' then
                  state_var1460 <= q_wait1180;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001")));
                  state_var1460 <= pause_getI1178;
                end if;
              when "1100" =>
                l := \$v1061\(0 to 31);
                \$v1188\ := \$arr963_ptr_take\;
                if \$v1188\(0) = '1' then
                  state_var1460 <= q_wait1187;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001")));
                  state_var1460 <= pause_getI1185;
                end if;
              when "1011" =>
                \$17_l\ := \$v1061\(0 to 31);
                \$v1195\ := \$arr963_ptr_take\;
                if \$v1195\(0) = '1' then
                  state_var1460 <= q_wait1194;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001")));
                  state_var1460 <= pause_getI1192;
                end if;
              when "0011" =>
                i := \$v1061\(0 to 31);
                \$v1203\ := \$arr963_ptr_take\;
                if \$v1203\(0) = '1' then
                  state_var1460 <= q_wait1202;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001")));
                  state_var1460 <= pause_getI1200;
                end if;
              when "0110" =>
                \$18_l\ := \$v1061\(0 to 31);
                \$v1208\ := \$arr963_ptr_take\;
                if \$v1208\(0) = '1' then
                  state_var1460 <= q_wait1207;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$v1204\ := \$18_l\ & vm_run_code247_arg(32 to 63);
                  \$arr963_ptr_write\ <= to_integer(unsigned(vm_run_code247_arg(0 to 31)));
                  \$arr963_write_request\ <= '1';
                  \$arr963_write\ <= "0100" & \$v1204\;
                  state_var1460 <= pause_setI1205;
                end if;
              when "1001" =>
                \$v1220\ := \$arr966_ptr_take\;
                if \$v1220\(0) = '1' then
                  state_var1460 <= q_wait1219;
                else
                  \$arr966_ptr_take\(0) := '1';
                  \$arr966_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(96 to 127) & "00000000000000000000000000000001")));
                  state_var1460 <= pause_getI1217;
                end if;
              when "0100" =>
                \$19_i\ := \$v1061\(0 to 31);
                \$v1228\ := \$arr962_ptr_take\;
                if \$v1228\(0) = '1' then
                  state_var1460 <= q_wait1227;
                else
                  \$arr962_ptr_take\(0) := '1';
                  \$arr962_ptr\ <= to_integer(unsigned(eclat_add(vm_run_code247_arg(32 to 63) & \$19_i\)));
                  state_var1460 <= pause_getI1225;
                end if;
              when "1010" =>
                \$20_l\ := \$v1061\(0 to 31);
                \$v752\ := vm_run_code247_arg(0 to 31) & vm_run_code247_arg(32 to 63) & eclat_sub(\$20_l\ & "00000000000000000000000000000001") & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
                \$v1060\ := ""&\$v752\(293);
                if \$v1060\(0) = '1' then
                  vm_run_code247_result := eclat_unit;
                  result1014 := vm_run_code247_result;
                  rdy1015 := eclat_true;
                  state_var1460 <= compute1016;
                else
                  vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                  state_var1460 <= vm_run_code247;
                end if;
              when "0111" =>
                \$v1240\ := eclat_eq(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & "00000000000000000000000000000000");
                if \$v1240\(0) = '1' then
                  \$v1239\ := \$arr963_ptr_take\;
                  if \$v1239\(0) = '1' then
                    state_var1460 <= q_wait1238;
                  else
                    \$arr963_ptr_take\(0) := '1';
                    \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001")));
                    state_var1460 <= pause_getI1236;
                  end if;
                else
                  \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
                  \$v1060\ := ""&\$v752\(293);
                  if \$v1060\(0) = '1' then
                    vm_run_code247_result := eclat_unit;
                    result1014 := vm_run_code247_result;
                    rdy1015 := eclat_true;
                    state_var1460 <= compute1016;
                  else
                    vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                    state_var1460 <= vm_run_code247;
                  end if;
                end if;
              when "0101" =>
                v := \$v1061\(0 to 67);
                \$v1244\ := \$arr963_ptr_take\;
                if \$v1244\(0) = '1' then
                  state_var1460 <= q_wait1243;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr_write\ <= to_integer(unsigned(vm_run_code247_arg(0 to 31)));
                  \$arr963_write_request\ <= '1';
                  \$arr963_write\ <= v;
                  state_var1460 <= pause_setI1241;
                end if;
              when "0010" =>
                \$21_i\ := \$v1061\(0 to 31);
                \$v1252\ := \$arr964_ptr_take\;
                if \$v1252\(0) = '1' then
                  state_var1460 <= q_wait1251;
                else
                  \$arr964_ptr_take\(0) := '1';
                  \$arr964_ptr\ <= to_integer(unsigned(\$21_i\));
                  state_var1460 <= pause_getI1249;
                end if;
              when "0001" =>
                \$22_i\ := \$v1061\(0 to 31);
                \$v1260\ := \$arr963_ptr_take\;
                if \$v1260\(0) = '1' then
                  state_var1460 <= q_wait1259;
                else
                  \$arr963_ptr_take\(0) := '1';
                  \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001")));
                  state_var1460 <= pause_getI1257;
                end if;
              when "0000" =>
                \$v752\ := vm_run_code247_arg(0 to 31) & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & eclat_add(vm_run_code247_arg(128 to 159) & "00000000000000000000000000000001") & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
                \$v1060\ := ""&\$v752\(293);
                if \$v1060\(0) = '1' then
                  vm_run_code247_result := eclat_unit;
                  result1014 := vm_run_code247_result;
                  rdy1015 := eclat_true;
                  state_var1460 <= compute1016;
                else
                  vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                  state_var1460 <= vm_run_code247;
                end if;
              when others =>
                eclat_print_string(of_string("Instr inconnu\n"));
                
                eclat_print_string(of_string("(exit) bye bye."));
                
                eclat_print_newline(eclat_unit);
                
                state_var1460 <= forever263939;
              end case;
            when pause_setI1017 =>
              \$arr962_write_request\ <= '0';
              state_var1460 <= pause_setII1018;
            when pause_setI1063 =>
              \$arr966_write_request\ <= '0';
              state_var1460 <= pause_setII1064;
            when pause_setI1067 =>
              \$arr966_write_request\ <= '0';
              state_var1460 <= pause_setII1068;
            when pause_setI1072 =>
              \$arr962_write_request\ <= '0';
              state_var1460 <= pause_setII1073;
            when pause_setI1077 =>
              \$arr963_write_request\ <= '0';
              state_var1460 <= pause_setII1078;
            when pause_setI1103 =>
              \$arr963_write_request\ <= '0';
              state_var1460 <= pause_setII1104;
            when pause_setI1122 =>
              \$arr963_write_request\ <= '0';
              state_var1460 <= pause_setII1123;
            when pause_setI1141 =>
              \$arr963_write_request\ <= '0';
              state_var1460 <= pause_setII1142;
            when pause_setI1153 =>
              \$arr963_write_request\ <= '0';
              state_var1460 <= pause_setII1154;
            when pause_setI1158 =>
              \$arr963_write_request\ <= '0';
              state_var1460 <= pause_setII1159;
            when pause_setI1170 =>
              \$arr963_write_request\ <= '0';
              state_var1460 <= pause_setII1171;
            when pause_setI1196 =>
              \$arr962_write_request\ <= '0';
              state_var1460 <= pause_setII1197;
            when pause_setI1205 =>
              \$arr963_write_request\ <= '0';
              state_var1460 <= pause_setII1206;
            when pause_setI1209 =>
              \$arr963_write_request\ <= '0';
              state_var1460 <= pause_setII1210;
            when pause_setI1221 =>
              \$arr963_write_request\ <= '0';
              state_var1460 <= pause_setII1222;
            when pause_setI1241 =>
              \$arr963_write_request\ <= '0';
              state_var1460 <= pause_setII1242;
            when pause_setI1245 =>
              \$arr963_write_request\ <= '0';
              state_var1460 <= pause_setII1246;
            when pause_setI1253 =>
              \$arr964_write_request\ <= '0';
              state_var1460 <= pause_setII1254;
            when pause_setII1018 =>
              \$arr962_ptr_take\(0) := '0';
              \$39_copy_args_to_heap257_arg\ := eclat_sub(\$39_copy_args_to_heap257_arg\(0 to 31) & "00000000000000000000000000000001") & \$39_copy_args_to_heap257_arg\(32 to 63) & eclat_add(\$39_copy_args_to_heap257_arg\(64 to 95) & "00000000000000000000000000000001") & \$39_copy_args_to_heap257_arg\(96 to 127) & \$39_copy_args_to_heap257_arg\(128 to 159);
              state_var1460 <= \$39_copy_args_to_heap257\;
            when pause_setII1064 =>
              \$arr966_ptr_take\(0) := '0';
              \$v752\ := eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001") & vm_run_code247_arg(160 to 191) & eclat_sub(\$v760\(0 to 31) & "00000000000000000000000000000001") & eclat_add(vm_run_code247_arg(96 to 127) & "00000000000000000000000000000001") & vm_run_code247_arg(128 to 159) & eclat_add(eclat_add(vm_run_code247_arg(160 to 191) & n) & "00000000000000000000000000000001") & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when pause_setII1068 =>
              \$arr966_ptr_take\(0) := '0';
              \$v1066\ := \$arr966_ptr_take\;
              if \$v1066\(0) = '1' then
                state_var1460 <= q_wait1065;
              else
                \$arr966_ptr_take\(0) := '1';
                \$arr966_ptr_write\ <= to_integer(unsigned(eclat_add(vm_run_code247_arg(96 to 127) & "00000000000000000000000000000001")));
                \$arr966_write_request\ <= '1';
                \$arr966_write\ <= eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001") & \$v760\(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127);
                state_var1460 <= pause_setI1063;
              end if;
            when pause_setII1073 =>
              \$arr962_ptr_take\(0) := '0';
              \$39_copy_args_to_heap257_arg\ := n & vm_run_code247_arg(0 to 31) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(0 to 31) & vm_run_code247_arg(32 to 63);
              state_var1460 <= \$39_copy_args_to_heap257\;
            when pause_setII1078 =>
              \$arr963_ptr_take\(0) := '0';
              \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & n) & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when pause_setII1104 =>
              \$arr963_ptr_take\(0) := '0';
              \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & n) & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when pause_setII1123 =>
              \$arr963_ptr_take\(0) := '0';
              \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & n) & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when pause_setII1142 =>
              \$arr963_ptr_take\(0) := '0';
              \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & n) & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when pause_setII1154 =>
              \$arr963_ptr_take\(0) := '0';
              \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & n) & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when pause_setII1159 =>
              \$arr963_ptr_take\(0) := '0';
              \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & n) & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when pause_setII1171 =>
              \$arr963_ptr_take\(0) := '0';
              \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & n) & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when pause_setII1197 =>
              \$arr962_ptr_take\(0) := '0';
              \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when pause_setII1206 =>
              \$arr963_ptr_take\(0) := '0';
              \$v752\ := eclat_add(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when pause_setII1210 =>
              \$arr963_ptr_take\(0) := '0';
              \$v752\ := eclat_add(\$v843\(0 to 31) & "00000000000000000000000000000001") & \$v843\(32 to 63) & \$v843\(64 to 95) & \$v843\(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when pause_setII1222 =>
              \$arr963_ptr_take\(0) := '0';
              \$v752\ := eclat_add(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when pause_setII1242 =>
              \$arr963_ptr_take\(0) := '0';
              \$v752\ := eclat_add(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when pause_setII1246 =>
              \$arr963_ptr_take\(0) := '0';
              \$v752\ := eclat_add(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when pause_setII1254 =>
              \$arr964_ptr_take\(0) := '0';
              \$v752\ := eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127) & vm_run_code247_arg(128 to 159) & vm_run_code247_arg(160 to 191) & vm_run_code247_arg(192 to 292) & ""&vm_run_code247_arg(293);
              \$v1060\ := ""&\$v752\(293);
              if \$v1060\(0) = '1' then
                vm_run_code247_result := eclat_unit;
                result1014 := vm_run_code247_result;
                rdy1015 := eclat_true;
                state_var1460 <= compute1016;
              else
                vm_run_code247_arg := \$v752\(0 to 31) & \$v752\(32 to 63) & eclat_add(\$v752\(64 to 95) & "00000000000000000000000000000001") & \$v752\(96 to 127) & \$v752\(128 to 159) & \$v752\(160 to 191) & \$v752\(192 to 292) & ""&\$v752\(293) & ""&vm_run_code247_arg(294);
                state_var1460 <= vm_run_code247;
              end if;
            when q_wait1019 =>
              \$v1020\ := \$arr962_ptr_take\;
              if \$v1020\(0) = '1' then
                state_var1460 <= q_wait1019;
              else
                \$arr962_ptr_take\(0) := '1';
                \$arr962_ptr_write\ <= to_integer(unsigned(\$39_copy_args_to_heap257_arg\(128 to 159)));
                \$arr962_write_request\ <= '1';
                \$arr962_write\ <= \$v13\;
                state_var1460 <= pause_setI1017;
              end if;
            when q_wait1023 =>
              \$v1024\ := \$arr963_ptr_take\;
              if \$v1024\(0) = '1' then
                state_var1460 <= q_wait1023;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$39_copy_args_to_heap257_arg\(96 to 127) & \$39_copy_args_to_heap257_arg\(0 to 31)) & "00000000000000000000000000000001")));
                state_var1460 <= pause_getI1021;
              end if;
            when q_wait1033 =>
              \$v1034\ := \$arr963_ptr_take\;
              if \$v1034\(0) = '1' then
                state_var1460 <= q_wait1033;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$41_div259_arg\(64 to 95) & "00000000000000000000000000000001") & \$41_div259_arg\(0 to 31))));
                state_var1460 <= pause_getI1031;
              end if;
            when q_wait1041 =>
              \$v1042\ := \$arr963_ptr_take\;
              if \$v1042\(0) = '1' then
                state_var1460 <= q_wait1041;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$42_mul260_arg\(64 to 95) & "00000000000000000000000000000001") & \$42_mul260_arg\(0 to 31))));
                state_var1460 <= pause_getI1039;
              end if;
            when q_wait1049 =>
              \$v1050\ := \$arr963_ptr_take\;
              if \$v1050\(0) = '1' then
                state_var1460 <= q_wait1049;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$43_sub261_arg\(64 to 95) & "00000000000000000000000000000001") & \$43_sub261_arg\(0 to 31))));
                state_var1460 <= pause_getI1047;
              end if;
            when q_wait1057 =>
              \$v1058\ := \$arr963_ptr_take\;
              if \$v1058\(0) = '1' then
                state_var1460 <= q_wait1057;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(\$44_add262_arg\(64 to 95) & "00000000000000000000000000000001") & \$44_add262_arg\(0 to 31))));
                state_var1460 <= pause_getI1055;
              end if;
            when q_wait1065 =>
              \$v1066\ := \$arr966_ptr_take\;
              if \$v1066\(0) = '1' then
                state_var1460 <= q_wait1065;
              else
                \$arr966_ptr_take\(0) := '1';
                \$arr966_ptr_write\ <= to_integer(unsigned(eclat_add(vm_run_code247_arg(96 to 127) & "00000000000000000000000000000001")));
                \$arr966_write_request\ <= '1';
                \$arr966_write\ <= eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001") & \$v760\(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127);
                state_var1460 <= pause_setI1063;
              end if;
            when q_wait1069 =>
              \$v1070\ := \$arr966_ptr_take\;
              if \$v1070\(0) = '1' then
                state_var1460 <= q_wait1069;
              else
                \$arr966_ptr_take\(0) := '1';
                \$arr966_ptr_write\ <= to_integer(unsigned(vm_run_code247_arg(96 to 127)));
                \$arr966_write_request\ <= '1';
                \$arr966_write\ <= eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001") & vm_run_code247_arg(32 to 63) & vm_run_code247_arg(64 to 95) & vm_run_code247_arg(96 to 127);
                state_var1460 <= pause_setI1067;
              end if;
            when q_wait1074 =>
              \$v1075\ := \$arr962_ptr_take\;
              if \$v1075\(0) = '1' then
                state_var1460 <= q_wait1074;
              else
                \$arr962_ptr_take\(0) := '1';
                \$v1071\ := vm_run_code247_arg(32 to 63);
                \$arr962_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_add(eclat_add(vm_run_code247_arg(160 to 191) & n) & "00000000000000000000000000000001") & "00000000000000000000000000000001")));
                \$arr962_write_request\ <= '1';
                \$arr962_write\ <= "0001" & \$v1071\&X"00000000";
                state_var1460 <= pause_setI1072;
              end if;
            when q_wait1079 =>
              \$v1080\ := \$arr963_ptr_take\;
              if \$v1080\(0) = '1' then
                state_var1460 <= q_wait1079;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001") & n)));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= "0000" & verif&"000"& X"000000000000000";
                state_var1460 <= pause_setI1077;
              end if;
            when q_wait1095 =>
              \$v1096\ := \$arr963_ptr_take\;
              if \$v1096\(0) = '1' then
                state_var1460 <= q_wait1095;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000011")));
                state_var1460 <= pause_getI1093;
              end if;
            when q_wait1099 =>
              \$v1100\ := \$arr963_ptr_take\;
              if \$v1100\(0) = '1' then
                state_var1460 <= q_wait1099;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000010")));
                state_var1460 <= pause_getI1097;
              end if;
            when q_wait1105 =>
              \$v1106\ := \$arr963_ptr_take\;
              if \$v1106\(0) = '1' then
                state_var1460 <= q_wait1105;
              else
                \$arr963_ptr_take\(0) := '1';
                \$v1102\ := eclat_gt(a & b);
                \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= "0000" & \$v1102\&"000"& X"000000000000000";
                state_var1460 <= pause_setI1103;
              end if;
            when q_wait1112 =>
              \$v1113\ := \$arr963_ptr_take\;
              if \$v1113\(0) = '1' then
                state_var1460 <= q_wait1112;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000010")));
                state_var1460 <= pause_getI1110;
              end if;
            when q_wait1119 =>
              \$v1120\ := \$arr963_ptr_take\;
              if \$v1120\(0) = '1' then
                state_var1460 <= q_wait1119;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000011")));
                state_var1460 <= pause_getI1117;
              end if;
            when q_wait1124 =>
              \$v1125\ := \$arr963_ptr_take\;
              if \$v1125\(0) = '1' then
                state_var1460 <= q_wait1124;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= "0001" & res&X"00000000";
                state_var1460 <= pause_setI1122;
              end if;
            when q_wait1131 =>
              \$v1132\ := \$arr963_ptr_take\;
              if \$v1132\(0) = '1' then
                state_var1460 <= q_wait1131;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000010")));
                state_var1460 <= pause_getI1129;
              end if;
            when q_wait1138 =>
              \$v1139\ := \$arr963_ptr_take\;
              if \$v1139\(0) = '1' then
                state_var1460 <= q_wait1138;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000011")));
                state_var1460 <= pause_getI1136;
              end if;
            when q_wait1143 =>
              \$v1144\ := \$arr963_ptr_take\;
              if \$v1144\(0) = '1' then
                state_var1460 <= q_wait1143;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= "0001" & res&X"00000000";
                state_var1460 <= pause_setI1141;
              end if;
            when q_wait1150 =>
              \$v1151\ := \$arr963_ptr_take\;
              if \$v1151\(0) = '1' then
                state_var1460 <= q_wait1150;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                state_var1460 <= pause_getI1148;
              end if;
            when q_wait1155 =>
              \$v1156\ := \$arr963_ptr_take\;
              if \$v1156\(0) = '1' then
                state_var1460 <= q_wait1155;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= "0001" & res&X"00000000";
                state_var1460 <= pause_setI1153;
              end if;
            when q_wait1160 =>
              \$v1161\ := \$arr963_ptr_take\;
              if \$v1161\(0) = '1' then
                state_var1460 <= q_wait1160;
              else
                \$arr963_ptr_take\(0) := '1';
                \$v1157\ := eclat_if(eclat_lt(resultat & "00000000000000000000000000000000") & eclat_mult(resultat & eclat_sub("00000000000000000000000000000000" & "00000000000000000000000000000001")) & resultat);
                \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= "0001" & \$v1157\&X"00000000";
                state_var1460 <= pause_setI1158;
              end if;
            when q_wait1167 =>
              \$v1168\ := \$arr963_ptr_take\;
              if \$v1168\(0) = '1' then
                state_var1460 <= q_wait1167;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                state_var1460 <= pause_getI1165;
              end if;
            when q_wait1172 =>
              \$v1173\ := \$arr963_ptr_take\;
              if \$v1173\(0) = '1' then
                state_var1460 <= q_wait1172;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr_write\ <= to_integer(unsigned(eclat_sub(eclat_sub(vm_run_code247_arg(0 to 31) & n) & "00000000000000000000000000000001")));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= "0001" & res&X"00000000";
                state_var1460 <= pause_setI1170;
              end if;
            when q_wait1180 =>
              \$v1181\ := \$arr963_ptr_take\;
              if \$v1181\(0) = '1' then
                state_var1460 <= q_wait1180;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001")));
                state_var1460 <= pause_getI1178;
              end if;
            when q_wait1187 =>
              \$v1188\ := \$arr963_ptr_take\;
              if \$v1188\(0) = '1' then
                state_var1460 <= q_wait1187;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001")));
                state_var1460 <= pause_getI1185;
              end if;
            when q_wait1194 =>
              \$v1195\ := \$arr963_ptr_take\;
              if \$v1195\(0) = '1' then
                state_var1460 <= q_wait1194;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001")));
                state_var1460 <= pause_getI1192;
              end if;
            when q_wait1198 =>
              \$v1199\ := \$arr962_ptr_take\;
              if \$v1199\(0) = '1' then
                state_var1460 <= q_wait1198;
              else
                \$arr962_ptr_take\(0) := '1';
                \$arr962_ptr_write\ <= to_integer(unsigned(eclat_add(vm_run_code247_arg(32 to 63) & i)));
                \$arr962_write_request\ <= '1';
                \$arr962_write\ <= var;
                state_var1460 <= pause_setI1196;
              end if;
            when q_wait1202 =>
              \$v1203\ := \$arr963_ptr_take\;
              if \$v1203\(0) = '1' then
                state_var1460 <= q_wait1202;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001")));
                state_var1460 <= pause_getI1200;
              end if;
            when q_wait1207 =>
              \$v1208\ := \$arr963_ptr_take\;
              if \$v1208\(0) = '1' then
                state_var1460 <= q_wait1207;
              else
                \$arr963_ptr_take\(0) := '1';
                \$v1204\ := \$18_l\ & vm_run_code247_arg(32 to 63);
                \$arr963_ptr_write\ <= to_integer(unsigned(vm_run_code247_arg(0 to 31)));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= "0100" & \$v1204\;
                state_var1460 <= pause_setI1205;
              end if;
            when q_wait1211 =>
              \$v1212\ := \$arr963_ptr_take\;
              if \$v1212\(0) = '1' then
                state_var1460 <= q_wait1211;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr_write\ <= to_integer(unsigned(\$v843\(0 to 31)));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= \$v151\;
                state_var1460 <= pause_setI1209;
              end if;
            when q_wait1215 =>
              \$v1216\ := \$arr963_ptr_take\;
              if \$v1216\(0) = '1' then
                state_var1460 <= q_wait1215;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001")));
                state_var1460 <= pause_getI1213;
              end if;
            when q_wait1219 =>
              \$v1220\ := \$arr966_ptr_take\;
              if \$v1220\(0) = '1' then
                state_var1460 <= q_wait1219;
              else
                \$arr966_ptr_take\(0) := '1';
                \$arr966_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(96 to 127) & "00000000000000000000000000000001")));
                state_var1460 <= pause_getI1217;
              end if;
            when q_wait1223 =>
              \$v1224\ := \$arr963_ptr_take\;
              if \$v1224\(0) = '1' then
                state_var1460 <= q_wait1223;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr_write\ <= to_integer(unsigned(vm_run_code247_arg(0 to 31)));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= temp;
                state_var1460 <= pause_setI1221;
              end if;
            when q_wait1227 =>
              \$v1228\ := \$arr962_ptr_take\;
              if \$v1228\(0) = '1' then
                state_var1460 <= q_wait1227;
              else
                \$arr962_ptr_take\(0) := '1';
                \$arr962_ptr\ <= to_integer(unsigned(eclat_add(vm_run_code247_arg(32 to 63) & \$19_i\)));
                state_var1460 <= pause_getI1225;
              end if;
            when q_wait1238 =>
              \$v1239\ := \$arr963_ptr_take\;
              if \$v1239\(0) = '1' then
                state_var1460 <= q_wait1238;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001")));
                state_var1460 <= pause_getI1236;
              end if;
            when q_wait1243 =>
              \$v1244\ := \$arr963_ptr_take\;
              if \$v1244\(0) = '1' then
                state_var1460 <= q_wait1243;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr_write\ <= to_integer(unsigned(vm_run_code247_arg(0 to 31)));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= v;
                state_var1460 <= pause_setI1241;
              end if;
            when q_wait1247 =>
              \$v1248\ := \$arr963_ptr_take\;
              if \$v1248\(0) = '1' then
                state_var1460 <= q_wait1247;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr_write\ <= to_integer(unsigned(vm_run_code247_arg(0 to 31)));
                \$arr963_write_request\ <= '1';
                \$arr963_write\ <= \$v170\;
                state_var1460 <= pause_setI1245;
              end if;
            when q_wait1251 =>
              \$v1252\ := \$arr964_ptr_take\;
              if \$v1252\(0) = '1' then
                state_var1460 <= q_wait1251;
              else
                \$arr964_ptr_take\(0) := '1';
                \$arr964_ptr\ <= to_integer(unsigned(\$21_i\));
                state_var1460 <= pause_getI1249;
              end if;
            when q_wait1255 =>
              \$v1256\ := \$arr964_ptr_take\;
              if \$v1256\(0) = '1' then
                state_var1460 <= q_wait1255;
              else
                \$arr964_ptr_take\(0) := '1';
                \$arr964_ptr_write\ <= to_integer(unsigned(\$22_i\));
                \$arr964_write_request\ <= '1';
                \$arr964_write\ <= \$v174\;
                state_var1460 <= pause_setI1253;
              end if;
            when q_wait1259 =>
              \$v1260\ := \$arr963_ptr_take\;
              if \$v1260\(0) = '1' then
                state_var1460 <= q_wait1259;
              else
                \$arr963_ptr_take\(0) := '1';
                \$arr963_ptr\ <= to_integer(unsigned(eclat_sub(vm_run_code247_arg(0 to 31) & "00000000000000000000000000000001")));
                state_var1460 <= pause_getI1257;
              end if;
            when q_wait1265 =>
              \$v1266\ := \$arr965_ptr_take\;
              if \$v1266\(0) = '1' then
                state_var1460 <= q_wait1265;
              else
                \$arr965_ptr_take\(0) := '1';
                \$arr965_ptr\ <= to_integer(unsigned(vm_run_code247_arg(64 to 95)));
                state_var1460 <= pause_getI1263;
              end if;
            when vm_run_code247 =>
              \$v1267\ := ""&vm_run_code247_arg(294);
              if \$v1267\(0) = '1' then
                eclat_print_string(of_string("[sp:"));
                
                eclat_print_int(vm_run_code247_arg(0 to 31));
                
                eclat_print_string(of_string("|env:"));
                
                eclat_print_int(vm_run_code247_arg(32 to 63));
                
                eclat_print_string(of_string("|pc:"));
                
                eclat_print_int(vm_run_code247_arg(64 to 95));
                
                eclat_print_string(of_string("|fp:"));
                
                eclat_print_int(vm_run_code247_arg(96 to 127));
                
                eclat_print_string(of_string("]"));
                
                eclat_print_string(of_string("|gp:"));
                
                eclat_print_int(vm_run_code247_arg(128 to 159));
                
                eclat_print_string(of_string("|hp:"));
                
                eclat_print_int(vm_run_code247_arg(128 to 159));
                
                eclat_print_newline(eclat_unit);
                
                \$v1266\ := \$arr965_ptr_take\;
                if \$v1266\(0) = '1' then
                  state_var1460 <= q_wait1265;
                else
                  \$arr965_ptr_take\(0) := '1';
                  \$arr965_ptr\ <= to_integer(unsigned(vm_run_code247_arg(64 to 95)));
                  state_var1460 <= pause_getI1263;
                end if;
              else
                \$v1266\ := \$arr965_ptr_take\;
                if \$v1266\(0) = '1' then
                  state_var1460 <= q_wait1265;
                else
                  \$arr965_ptr_take\(0) := '1';
                  \$arr965_ptr\ <= to_integer(unsigned(vm_run_code247_arg(64 to 95)));
                  state_var1460 <= pause_getI1263;
                end if;
              end if;
            when compute1016 =>
              rdy1015 := eclat_false;
              eclat_print_string(of_string("START (cy="));
              
              eclat_print_int(cy);
              
              eclat_print_string(of_string(")"));
              
              eclat_print_newline(eclat_unit);
              
              \$v1268\ := eclat_unit;
              vm_run_code247_arg := "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & "00000000000000000000000000000000" & eclat_false & "00000000000000000000000000000000" & "0010" & \$v1268\&"000"& X"000000000000000" & eclat_false & argument;
              state_var1460 <= vm_run_code247;
            end case;
            \$v1270\ := eclat_not(rdy1015);
            if \$v1270\(0) = '1' then
              result1014 := eclat_unit;
            end if;
            \$v711\ := result1014 & rdy1015;
            \$v1013\ := ""&\$v711\(1);
            if \$v1013\(0) = '1' then
              eclat_print_string(of_string("END (cy="));
              
              eclat_print_int(cy);
              
              eclat_print_string(of_string(")"));
              
              eclat_print_newline(eclat_unit);
              
              result967 := eclat_unit;
              eclat_print_newline(eclat_unit);
              
              rdy968 := eclat_true;
              \state\ <= compute969;
            else
              result967 := eclat_unit;
              rdy968 := eclat_true;
              \state\ <= compute969;
            end if;
          end case;
          
          result <= result967;
          rdy <= rdy968;
          
        end if;
      end if;
    end if;
  end process;
end architecture;
